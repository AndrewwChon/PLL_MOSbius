** sch_path: /foss/designs/libs/xp_core_analog/xp_programmable_basic_pump_flatten/xp_programmable_basic_pump.sch
.subckt xp_programmable_basic_pump VDD VSS up down iref out s3 s4 s1 s2
*.PININFO VDD:B VSS:B up:B down:B iref:B out:B s3:B s4:B s1:B s2:B
M6 out net5 net4 VSS nfet_03v3 L=0.5u W=14.0u nf=2 m=1
M8 net7 upb VDD VDD pfet_03v3 L=0.5u W=42.0u nf=6 m=1
M10 net6 VSS VDD VDD pfet_03v3 L=0.5u W=42.0u nf=6 m=1
x1 up VDD upb VSS inv1u05u
x2 net3 VSS s1 net8 s1b VDD pass1u05u
x4 iref VSS s1 net5 s1b VDD pass1u05u
x6 s1 VDD s1b VSS inv1u05u
x7 s2 VDD s2b VSS inv1u05u
x8 s3 VDD s3b VSS inv1u05u
x9 s4 VDD s4b VSS inv1u05u
M12 out net10 net9 VSS nfet_03v3 L=0.5u W=14.0u nf=2 m=2
M14 net11 upb VDD VDD pfet_03v3 L=0.5u W=42.0u nf=6 m=2
x12 net3 VSS s2 net12 s2b VDD pass1u05u
x14 iref VSS s2 net10 s2b VDD pass1u05u
M16 out net14 net13 VSS nfet_03v3 L=0.5u W=14.0u nf=2 m=4
M18 net15 upb VDD VDD pfet_03v3 L=0.5u W=42.0u nf=6 m=4
x16 net3 VSS s3 net16 s3b VDD pass1u05u
x18 iref VSS s3 net14 s3b VDD pass1u05u
M19 out net20 net19 VDD pfet_03v3 L=0.5u W=42.0u nf=6 m=8
M20 out net18 net17 VSS nfet_03v3 L=0.5u W=14.0u nf=2 m=8
M22 net19 upb VDD VDD pfet_03v3 L=0.5u W=42.0u nf=6 m=8
x20 net3 VSS s4 net20 s4b VDD pass1u05u
x22 iref VSS s4 net18 s4b VDD pass1u05u
M2 iref iref net1 VSS nfet_03v3 L=0.5u W=14.0u nf=2 m=1
M9 net3 net3 net6 VDD pfet_03v3 L=0.5u W=42.0u nf=6 m=1
M1 out net8 net7 VDD pfet_03v3 L=0.5u W=42.0u nf=6 m=1
M11 out net12 net11 VDD pfet_03v3 L=0.5u W=42.0u nf=6 m=2
M15 out net16 net15 VDD pfet_03v3 L=0.5u W=42.0u nf=6 m=4
M3 net1 VDD VSS VSS nfet_03v3 L=0.5u W=14.0u nf=2 m=1
M4 net2 VDD VSS VSS nfet_03v3 L=0.5u W=14.0u nf=2 m=1
M5 net3 iref net2 VSS nfet_03v3 L=0.5u W=14.0u nf=2 m=1
M21 net4 down VSS VSS nfet_03v3 L=0.5u W=14.0u nf=2 m=1
M7 net9 down VSS VSS nfet_03v3 L=0.5u W=14.0u nf=2 m=2
M13 net13 down VSS VSS nfet_03v3 L=0.5u W=14.0u nf=2 m=4
M17 net17 down VSS VSS nfet_03v3 L=0.5u W=14.0u nf=2 m=8
M23 VSS VSS VSS VSS nfet_03v3 L=0.5u W=14.0u nf=2 m=6
M24 VSS VSS VSS VSS nfet_03v3 L=0.5u W=14.0u nf=2 m=6
M26 net5 s1b VSS VSS nfet_03v3 L=0.5u W=1.0u nf=1 m=1
M29 net8 s1 VDD VDD pfet_03v3 L=0.5u W=1.0u nf=1 m=1
M33 VDD VDD VDD VDD pfet_03v3 L=0.5u W=42.0u nf=6 m=4
M34 VDD VDD VDD VDD pfet_03v3 L=0.5u W=7.0u nf=1 m=6
M36 VDD VDD VDD VDD pfet_03v3 L=0.5u W=7.0u nf=1 m=6
M25 net10 s2b VSS VSS nfet_03v3 L=0.5u W=1.0u nf=1 m=1
M27 net14 s3b VSS VSS nfet_03v3 L=0.5u W=1.0u nf=1 m=1
M28 net18 s4b VSS VSS nfet_03v3 L=0.5u W=1.0u nf=1 m=1
M30 net12 s2 VDD VDD pfet_03v3 L=0.5u W=1.0u nf=1 m=1
M31 net16 s3 VDD VDD pfet_03v3 L=0.5u W=1.0u nf=1 m=1
M32 net20 s4 VDD VDD pfet_03v3 L=0.5u W=1.0u nf=1 m=1
.ends

* expanding   symbol:  libs/core_analog/inv1u05u/inv1u05u.sym # of pins=4
** sym_path: /foss/designs/libs/core_analog/inv1u05u/inv1u05u.sym
** sch_path: /foss/designs/libs/core_analog/inv1u05u/inv1u05u.sch
.subckt inv1u05u in vdd out vss
*.PININFO in:B out:B vss:B vdd:B
M1 out in vdd vdd pfet_03v3 L=0.5u W=3.0u nf=1 m=1
M2 out in vss vss nfet_03v3 L=0.5u W=1.0u nf=1 m=1
.ends


* expanding   symbol:  libs/core_analog/pass1u05u/pass1u05u.sym # of pins=6
** sym_path: /foss/designs/libs/core_analog/pass1u05u/pass1u05u.sym
** sch_path: /foss/designs/libs/core_analog/pass1u05u/pass1u05u.sch
.subckt pass1u05u ind vss clkn ins clkp vdd
*.PININFO ind:B ins:B clkn:B clkp:B vdd:B vss:B
M1 ind clkp ins vdd pfet_03v3 L=0.5u W=3.0u nf=1 m=1
M2 ind clkn ins vss nfet_03v3 L=0.5u W=1.0u nf=1 m=1
.ends

