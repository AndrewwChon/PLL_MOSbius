* NGSPICE file created from top_level_20250912_sc.ext - technology: gf180mcuD

.subckt nfet$280 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$258 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$261 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$278 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt nfet$276 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$259 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$257 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$260 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$279 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$277 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt asc_drive_buffer_up vss out in vdd
Xnfet$280_0 in vss m1_n566_1318# vss nfet$280
Xpfet$258_0 m1_778_712# vdd vdd m1_778_712# m1_506_712# m1_506_712# m1_778_712# vdd
+ m1_506_712# m1_506_712# pfet$258
Xpfet$261_0 vdd vdd m1_n566_1318# in pfet$261
Xnfet$278_0 m1_n30_1318# vss m1_506_712# vss nfet$278
Xnfet$276_0 m1_778_712# vss m1_506_712# m1_506_712# m1_506_712# m1_778_712# m1_778_712#
+ vss m1_506_712# vss nfet$276
Xpfet$259_0 vdd vdd m1_506_712# m1_n30_1318# pfet$259
Xpfet$257_0 out out m1_778_712# vdd m1_778_712# out vdd vdd m1_778_712# out m1_778_712#
+ m1_778_712# out m1_778_712# vdd m1_778_712# vdd m1_778_712# pfet$257
Xpfet$260_0 vdd vdd m1_n30_1318# m1_n566_1318# pfet$260
Xnfet$279_0 m1_n566_1318# vss m1_n30_1318# vss nfet$279
Xnfet$277_0 out out vss m1_778_712# m1_778_712# out vss m1_778_712# m1_778_712# m1_778_712#
+ out m1_778_712# m1_778_712# out vss m1_778_712# vss vss nfet$277
.ends

.subckt pfet$196 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$238 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$212 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$224 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$217 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$231 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$207 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$214 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$215 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$221 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$197 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$213 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$220 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$205 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$202 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$211 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$199 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$243 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$228 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$210 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$236 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$203 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$229 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$241 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$226 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$234 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$219 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$201 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$227 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$224 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$232 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$217 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$200 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$225 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$218 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$222 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$230 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$215 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$223 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$208 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$216 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$220 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$246 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$213 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$239 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$221 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$206 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$198 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$214 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$244 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$219 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$211 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$237 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$204 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$242 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$227 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$235 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$228 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$225 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$240 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$233 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$218 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$226 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$223 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$216 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$209 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$247 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$222 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$245 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$212 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt asc_dual_psd_def_20250809 vdd vss pd1 pd2 pd3 pd4 pd5 pd6 pd7 pd8 pd9 fout
+ sd1 sd2 sd3 sd4 sd5 sd6 sd7 sd8 sd9 fin define
Xpfet$196_7 vdd vdd m1_7232_25662# m1_7095_25858# pfet$196
Xnfet$238_1 m1_n1927_20274# m1_n1927_20274# vss vss m1_n2445_20470# vss nfet$238
Xnfet$212_72 m1_23827_25858# m1_25912_25658# m1_26705_24542# vss nfet$212
Xnfet$212_61 m1_23964_25662# m1_24808_24224# m1_25912_25658# vss nfet$212
Xnfet$212_50 m1_n7513_20152# vss m1_21241_24346# vss nfet$212
Xnfet$224_7 m1_488_21786# m1_488_21786# vss vss m1_n674_21586# vss nfet$224
Xnfet$217_6 m1_9015_17714# vss m1_12935_19550# vss nfet$217
Xnfet$231_8 m1_3015_15778# m1_3015_15778# m1_2905_18030# m1_2905_18030# m1_3141_17358#
+ vss nfet$231
Xnfet$217_17 m1_21880_15478# vss m1_25722_20152# vss nfet$217
Xpfet$196_49 vdd m1_20126_25858# vdd m1_21729_25658# pfet$196
Xpfet$196_38 vdd vdd m1_16085_25662# m1_15943_25858# pfet$196
Xpfet$196_27 vdd vdd m1_11278_25858# m1_7522_21786# pfet$196
Xpfet$196_16 vdd vdd m1_5771_21786# pd3 pfet$196
Xpfet$207_4 vdd m1_34093_19792# vdd m1_32818_20470# pfet$207
Xpfet$214_5 vdd m1_26217_17714# vdd m1_27292_16202# pfet$214
Xnfet$215_3 m1_n7513_20152# vss m1_9944_16080# vss nfet$215
Xpfet$221_6 vdd vdd m1_n6973_21481# m1_n6839_21786# pfet$221
Xpfet$197_92 vdd m1_15454_18030# vdd m1_14127_16080# pfet$197
Xpfet$197_81 vdd vdd m1_13668_17714# m1_14127_16080# pfet$197
Xpfet$197_70 vdd vdd m1_18824_17836# m1_18665_17343# pfet$197
Xnfet$213_0 m1_n1133_21590# m1_n1133_21590# m1_354_22513# m1_354_22513# m1_n674_21586#
+ vss nfet$213
Xnfet$220_1 m1_n789_25858# vss m1_n647_25662# vss nfet$220
Xpfet$205_1 vdd m1_n789_25858# vdd m1_814_25658# pfet$205
Xpfet$202_13 vdd vdd m1_16452_19550# m1_13198_17714# pfet$202
Xpfet$197_103 vdd m1_14743_16202# m1_14258_17518# m1_14641_17836# pfet$197
Xnfet$215_72 m1_17851_17714# vss m1_18441_17518# vss nfet$215
Xnfet$215_61 m1_20104_16080# vss m1_19747_15778# vss nfet$215
Xnfet$215_50 m1_25747_17714# vss m1_22848_17343# vss nfet$215
Xnfet$211_19 m1_21729_25658# m1_21729_25658# vss vss m1_22188_25502# vss nfet$211
Xpfet$199_27 vdd vdd vdd m1_20407_19850# m1_22205_20152# m1_22205_20152# pfet$199
Xpfet$199_16 vdd vdd vdd m1_28077_19550# m1_26063_15478# m1_26063_15478# pfet$199
Xpfet$196_8 vdd vdd m1_8076_24224# m1_7456_23922# pfet$196
Xnfet$238_2 m1_n3206_20274# m1_n3206_20274# vss vss m1_n3724_20470# vss nfet$238
Xnfet$212_73 m1_24309_25858# vss m1_21590_21786# vss nfet$212
Xnfet$212_62 m1_24188_23922# vss m1_24808_24224# vss nfet$212
Xnfet$212_51 m1_19644_25858# m1_21729_25658# m1_22522_24542# vss nfet$212
Xnfet$212_40 m1_15598_25662# m1_16442_24224# m1_17546_25658# vss nfet$212
Xnfet$224_8 m1_25739_21786# m1_25739_21786# vss vss m1_24577_21586# vss nfet$224
Xnfet$217_7 m1_5148_15478# vss m1_11654_20152# vss nfet$217
Xnfet$231_9 m1_2194_16202# m1_2194_16202# vss vss m1_1676_16398# vss nfet$231
Xpfet$196_39 vdd vdd m1_15598_25662# m1_15461_25858# pfet$196
Xpfet$196_28 vdd m1_11639_23922# m1_11903_24542# m1_11278_25858# pfet$196
Xpfet$196_17 vdd vdd m1_7577_25858# m1_8692_24346# pfet$196
Xnfet$243_0 m1_n8283_20611# vss m1_n8283_19850# vss nfet$243
Xpfet$228_0 vdd vdd m1_n8145_21908# m1_n6839_20152# pfet$228
Xpfet$214_6 vdd vdd m1_28003_18030# m1_28113_15778# pfet$214
Xpfet$207_5 vdd vdd m1_34093_19792# m1_32818_21586# pfet$207
Xnfet$215_4 m1_10299_17343# m1_10560_16202# m1_10075_17518# vss nfet$215
Xpfet$221_7 vdd vdd m1_n6839_21786# m1_n6380_21786# pfet$221
Xpfet$197_93 vdd m1_23820_18030# vdd m1_22493_16080# pfet$197
Xpfet$197_82 vdd m1_13668_17714# vdd m1_14743_16202# pfet$197
Xpfet$197_71 vdd vdd m1_19747_15778# m1_20104_16080# pfet$197
Xpfet$197_60 vdd vdd m1_n194_15778# m1_n3064_17714# pfet$197
Xnfet$213_1 m1_n1263_21786# m1_n1263_21786# m1_354_22513# m1_354_22513# m1_n42_21586#
+ vss nfet$213
Xnfet$220_2 m1_n1271_25858# vss m1_n1134_25662# vss nfet$220
Xpfet$205_2 vdd vdd m1_n789_25858# m1_326_24346# pfet$205
Xpfet$202_14 vdd vdd m1_23486_19550# m1_21564_17714# pfet$202
Xpfet$197_104 vdd vdd m1_14127_16080# m1_n7513_20152# pfet$197
Xpfet$210_0 vdd m1_34093_22102# vdd m1_28490_22513# pfet$210
Xnfet$215_73 m1_13668_17714# vss m1_16538_15778# vss nfet$215
Xnfet$215_62 m1_18665_17343# m1_20721_15778# m1_20104_16080# vss nfet$215
Xnfet$215_51 m1_n7513_20152# vss m1_22493_16080# vss nfet$215
Xnfet$215_40 m1_n2250_17343# m1_n194_15778# m1_n811_16080# vss nfet$215
Xpfet$199_28 vdd vdd vdd m1_21043_19550# m1_17697_15478# m1_17697_15478# pfet$199
Xpfet$199_17 vdd m1_n3822_20130# m1_n3822_20130# m1_28077_19550# m1_25747_17714# m1_25747_17714#
+ pfet$199
Xnfet$238_3 m1_n6973_21481# m1_n6973_21481# m1_n6839_20152# m1_n6839_20152# m1_n6282_20470#
+ vss nfet$238
Xpfet$196_9 vdd m1_7719_25662# m1_7456_23922# m1_7232_25662# pfet$196
Xnfet$212_74 pd8 vss m1_23356_21786# vss nfet$212
Xnfet$212_63 m1_14556_21786# vss m1_19644_25858# vss nfet$212
Xnfet$212_52 m1_20126_25858# vss m1_22522_24542# vss nfet$212
Xnfet$212_41 pd5 vss m1_12805_21786# vss nfet$212
Xnfet$212_30 m1_n7513_20152# vss m1_17058_24346# vss nfet$212
Xnfet$224_9 m1_25107_21786# m1_25107_21786# vss vss m1_23945_21586# vss nfet$224
Xnfet$217_8 m1_n7383_17599# vss m1_n1133_19550# vss nfet$217
Xpfet$196_29 vdd vdd m1_11903_24542# m1_12259_24224# pfet$196
Xpfet$196_18 vdd vdd m1_11415_25662# m1_11278_25858# pfet$196
Xnfet$243_1 m1_n7513_20152# m1_n8283_19850# vss vss nfet$243
Xnfet$236_0 m1_n10452_25858# m1_n10452_25858# m1_n7186_25858# m1_n7186_25858# m1_n6629_25502#
+ vss nfet$236
Xnfet$215_5 m1_10458_17836# m1_11738_16080# m1_11271_18030# vss nfet$215
Xpfet$214_7 vdd m1_28003_18030# vdd m1_26676_16080# pfet$214
Xpfet$207_6 vdd vdd m1_31535_19792# m1_14422_22513# pfet$207
Xpfet$197_94 vdd vdd m1_22624_17518# m1_22034_17714# pfet$197
Xpfet$197_83 vdd m1_16538_15778# m1_15921_16080# m1_14641_17836# pfet$197
Xpfet$197_72 vdd m1_20721_15778# m1_20104_16080# m1_18824_17836# pfet$197
Xpfet$197_61 vdd m1_n811_16080# m1_n1278_18030# m1_n2250_17343# pfet$197
Xpfet$197_50 vdd m1_n1168_15778# m1_n1989_16202# m1_n2250_17343# pfet$197
Xpfet$205_3 vdd m1_n646_24542# vdd m1_326_24346# pfet$205
Xnfet$213_2 m1_9288_21786# m1_9288_21786# m1_9645_21447# m1_9645_21447# m1_10509_21586#
+ vss nfet$213
Xnfet$220_3 m1_n7513_20152# vss m1_326_24346# vss nfet$220
Xpfet$202_15 vdd vdd m1_22205_20152# m1_17697_15478# pfet$202
Xpfet$197_105 vdd vdd m1_14258_17518# m1_13668_17714# pfet$197
Xpfet$210_1 vdd vdd m1_34093_22102# m1_34843_21786# pfet$210
Xnfet$215_74 m1_14482_17343# vss m1_14641_17836# vss nfet$215
Xnfet$215_63 m1_13668_17714# vss m1_14258_17518# vss nfet$215
Xnfet$215_52 m1_23007_17836# m1_24287_16080# m1_23820_18030# vss nfet$215
Xnfet$215_30 sd6 vss m1_5148_15478# vss nfet$215
Xnfet$215_41 m1_n2091_17836# m1_n1168_15778# m1_n1989_16202# vss nfet$215
Xpfet$203_0 vdd vdd m1_n7401_15478# sd9 pfet$203
Xpfet$199_29 vdd vdd vdd m1_23924_19850# m1_25722_20152# m1_25722_20152# pfet$199
Xpfet$199_18 vdd vdd vdd m1_27441_19850# m1_29239_20152# m1_29239_20152# pfet$199
Xnfet$238_4 m1_2590_19404# m1_2590_19404# vss vss m1_n2445_21430# vss nfet$238
Xnfet$212_75 m1_28371_23922# vss m1_28991_24224# vss nfet$212
Xnfet$212_64 m1_19644_25858# vss m1_19781_25662# vss nfet$212
Xnfet$212_53 m1_23827_25858# m1_24451_25662# m1_24188_23922# vss nfet$212
Xnfet$212_42 m1_15943_25858# vss m1_16085_25662# vss nfet$212
Xnfet$212_31 m1_15943_25858# vss m1_18339_24542# vss nfet$212
Xnfet$217_9 m1_25747_17714# vss m1_27003_19550# vss nfet$217
Xnfet$212_20 pd3 vss m1_5771_21786# vss nfet$212
Xnfet$229_0 m1_34093_22102# vss fout vss nfet$229
Xnfet$243_2 m1_n8145_21908# vss m1_n8283_20611# vss nfet$243
Xnfet$236_1 m1_n6111_25858# m1_n6111_25858# vss vss m1_n6629_25502# vss nfet$236
Xpfet$196_19 vdd vdd m1_7095_25858# m1_4005_21786# pfet$196
Xnfet$215_6 m1_6116_17343# vss m1_6275_17836# vss nfet$215
Xpfet$207_7 vdd vdd m1_31535_22102# m1_354_22513# pfet$207
Xpfet$197_95 vdd vdd m1_21564_17714# m1_22034_17714# pfet$197
Xpfet$197_84 vdd vdd m1_17381_17714# m1_17851_17714# pfet$197
Xpfet$197_73 vdd vdd m1_16538_15778# m1_13668_17714# pfet$197
Xpfet$197_62 vdd vdd m1_23007_17836# m1_22848_17343# pfet$197
Xpfet$197_40 vdd m1_10560_16202# m1_10075_17518# m1_10458_17836# pfet$197
Xpfet$197_51 vdd vdd m1_n1168_15778# m1_n811_16080# pfet$197
Xnfet$213_3 m1_9418_21590# m1_9418_21590# m1_9645_21447# m1_9645_21447# m1_9877_21586#
+ vss nfet$213
Xnfet$220_4 m1_n789_25858# vss m1_1607_24542# vss nfet$220
Xpfet$205_4 vdd vdd m1_32675_25947# m1_33790_24346# pfet$205
Xpfet$197_106 vdd vdd m1_14482_17343# m1_17381_17714# pfet$197
Xpfet$202_16 vdd vdd m1_19969_19550# m1_17381_17714# pfet$202
Xnfet$211_0 m1_4509_24346# m1_4509_24346# vss vss m1_3991_24542# vss nfet$211
Xpfet$210_2 vdd vdd m1_30256_22102# m1_7388_22513# pfet$210
Xpfet$203_1 vdd vdd m1_21880_15478# sd2 pfet$203
Xnfet$215_31 m1_1933_17343# m1_3989_15778# m1_3372_16080# vss nfet$215
Xnfet$215_20 m1_1119_17714# vss m1_1709_17518# vss nfet$215
Xnfet$215_42 m1_n811_16080# vss m1_n1168_15778# vss nfet$215
Xnfet$215_75 sd3 vss m1_17697_15478# vss nfet$215
Xnfet$215_64 m1_13668_17714# vss m1_13198_17714# vss nfet$215
Xnfet$215_53 m1_22848_17343# vss m1_23007_17836# vss nfet$215
Xpfet$199_19 vdd m1_n3822_20130# m1_n3822_20130# m1_27441_19850# m1_27003_19550# m1_27003_19550#
+ pfet$199
Xnfet$238_5 m1_6107_19404# m1_6107_19404# m1_n5227_21418# m1_n5227_21418# m1_n2445_21430#
+ vss nfet$238
Xnfet$212_76 m1_28492_25858# vss m1_28634_25662# vss nfet$212
Xnfet$212_65 m1_28492_25858# vss m1_25107_21786# vss nfet$212
Xnfet$212_54 m1_24309_25858# vss m1_24451_25662# vss nfet$212
Xnfet$212_43 m1_15461_25858# vss m1_15598_25662# vss nfet$212
Xnfet$212_32 m1_15461_25858# m1_17546_25658# m1_18339_24542# vss nfet$212
Xnfet$212_21 m1_11278_25858# m1_11902_25662# m1_11639_23922# vss nfet$212
Xnfet$212_10 m1_7577_25858# vss m1_9973_24542# vss nfet$212
Xnfet$243_3 m1_n8283_19850# m1_n8283_20611# vss vss nfet$243
Xnfet$215_7 m1_9485_17714# vss m1_10075_17518# vss nfet$215
Xnfet$241_0 m1_n10933_25858# m1_n8848_25658# m1_n8055_24542# vss nfet$241
Xpfet$197_96 vdd vdd m1_18665_17343# m1_21564_17714# pfet$197
Xpfet$197_85 vdd m1_18926_16202# m1_18441_17518# m1_18824_17836# pfet$197
Xpfet$197_74 vdd vdd m1_14641_17836# m1_14482_17343# pfet$197
Xpfet$197_63 vdd m1_23930_15778# m1_23109_16202# m1_22848_17343# pfet$197
Xpfet$197_30 vdd vdd m1_1933_17343# m1_4832_17714# pfet$197
Xpfet$197_41 vdd vdd m1_10075_17518# m1_9485_17714# pfet$197
Xpfet$197_52 vdd m1_n3064_17714# vdd m1_n1989_16202# pfet$197
Xpfet$226_0 vdd vdd m1_n5227_20152# m1_n2543_20130# pfet$226
Xnfet$213_4 m1_5901_21590# m1_5901_21590# m1_7388_22513# m1_7388_22513# m1_6360_21586#
+ vss nfet$213
Xnfet$220_5 m1_n789_25858# vss m1_488_21786# vss nfet$220
Xpfet$205_5 vdd m1_32675_25947# vdd m1_34278_25658# pfet$205
Xnfet$220_10 m1_32675_25947# vss m1_35071_24542# vss nfet$220
Xpfet$202_17 vdd vdd m1_25722_20152# m1_21880_15478# pfet$202
Xpfet$197_107 vdd m1_15921_16080# m1_15454_18030# m1_14482_17343# pfet$197
Xpfet$203_2 vdd vdd m1_26063_15478# sd1 pfet$203
Xpfet$210_3 vdd m1_31535_22102# vdd m1_3871_22513# pfet$210
Xnfet$211_1 m1_3893_24224# m1_3893_24224# m1_3537_24542# m1_3537_24542# m1_3991_24542#
+ vss nfet$211
Xnfet$215_76 m1_14482_17343# m1_16538_15778# m1_15921_16080# vss nfet$215
Xnfet$215_65 m1_14482_17343# m1_14743_16202# m1_14258_17518# vss nfet$215
Xnfet$231_20 m1_22493_16080# m1_22493_16080# m1_22034_17714# m1_22034_17714# m1_22591_16398#
+ vss nfet$231
Xnfet$215_54 m1_22848_17343# m1_23109_16202# m1_22624_17518# vss nfet$215
Xnfet$215_32 m1_2092_17836# m1_3015_15778# m1_2194_16202# vss nfet$215
Xnfet$215_21 m1_1933_17343# m1_2194_16202# m1_1709_17518# vss nfet$215
Xnfet$215_10 m1_11738_16080# vss m1_11381_15778# vss nfet$215
Xnfet$215_43 sd8 vss m1_n3218_15478# vss nfet$215
Xnfet$238_6 m1_n5764_21786# m1_n5764_21786# vss vss m1_n6282_21430# vss nfet$238
Xnfet$212_77 m1_28010_25858# vss m1_28147_25662# vss nfet$212
Xnfet$212_66 m1_28010_25858# m1_30095_25658# m1_30888_24542# vss nfet$212
Xnfet$212_55 m1_23827_25858# vss m1_23964_25662# vss nfet$212
Xnfet$212_44 m1_15822_23922# vss m1_16442_24224# vss nfet$212
Xnfet$212_33 m1_11760_25858# vss m1_14156_24542# vss nfet$212
Xnfet$212_22 m1_11760_25858# vss m1_11902_25662# vss nfet$212
Xnfet$212_11 m1_7522_21786# vss m1_11278_25858# vss nfet$212
Xnfet$215_8 m1_7555_16080# vss m1_7198_15778# vss nfet$215
Xnfet$234_0 m1_n6274_17836# m1_n4994_16080# m1_n5461_18030# vss nfet$234
Xnfet$241_1 m1_n10796_25662# m1_n10572_23922# m1_n10308_24542# vss nfet$241
Xpfet$197_20 vdd vdd m1_1119_17714# m1_1578_16080# pfet$197
Xpfet$226_1 vdd m1_n4485_20152# vdd m1_n3206_20274# pfet$226
Xpfet$219_0 vdd vdd m1_n7320_25516# m1_n7186_25858# pfet$219
Xpfet$197_97 vdd vdd m1_22493_16080# m1_n7513_20152# pfet$197
Xpfet$197_86 vdd m1_19637_18030# vdd m1_18310_16080# pfet$197
Xpfet$197_75 vdd vdd m1_17697_15478# sd3 pfet$197
Xpfet$197_64 vdd vdd m1_23930_15778# m1_24287_16080# pfet$197
Xnfet$220_6 m1_n910_23922# vss m1_n290_24224# vss nfet$220
Xpfet$197_31 vdd m1_3372_16080# m1_2905_18030# m1_1933_17343# pfet$197
Xpfet$197_42 vdd m1_11271_18030# vdd m1_9944_16080# pfet$197
Xpfet$197_53 vdd vdd m1_n3218_15478# sd8 pfet$197
Xnfet$213_5 m1_2254_21786# m1_2254_21786# m1_3871_22513# m1_3871_22513# m1_3475_21586#
+ vss nfet$213
Xpfet$205_6 vdd vdd m1_32818_24542# m1_33174_24224# pfet$205
Xnfet$220_11 m1_32554_23922# vss m1_33174_24224# vss nfet$220
Xpfet$210_4 vdd m1_30256_22102# vdd m1_9645_21447# pfet$210
Xpfet$197_108 vdd vdd m1_15454_18030# m1_15564_15778# pfet$197
Xnfet$211_2 m1_4997_25658# m1_4997_25658# vss vss m1_5456_25502# vss nfet$211
Xnfet$215_77 sd4 vss m1_13514_15478# vss nfet$215
Xnfet$215_66 m1_n7513_20152# vss m1_14127_16080# vss nfet$215
Xnfet$231_21 m1_14127_16080# m1_14127_16080# vss vss m1_15690_17358# vss nfet$231
Xnfet$215_55 m1_22034_17714# vss m1_24904_15778# vss nfet$215
Xnfet$215_44 m1_n2091_17836# m1_n811_16080# m1_n1278_18030# vss nfet$215
Xnfet$215_33 sd7 vss m1_965_15478# vss nfet$215
Xnfet$231_10 m1_1578_16080# m1_1578_16080# m1_1119_17714# m1_1119_17714# m1_1676_16398#
+ vss nfet$231
Xnfet$215_22 m1_6116_17343# m1_6377_16202# m1_5892_17518# vss nfet$215
Xnfet$215_11 m1_10299_17343# m1_12355_15778# m1_11738_16080# vss nfet$215
Xpfet$201_0 vdd vdd m1_n6274_17836# m1_n6433_17343# pfet$201
Xnfet$238_7 m1_n3822_21786# m1_n3822_21786# m1_n4485_21904# m1_n4485_21904# m1_n3724_21430#
+ vss nfet$238
Xnfet$212_12 m1_7577_25858# vss m1_7522_21786# vss nfet$212
Xnfet$212_78 m1_28010_25858# m1_28634_25662# m1_28371_23922# vss nfet$212
Xnfet$212_67 m1_28492_25858# vss m1_30888_24542# vss nfet$212
Xnfet$212_56 m1_19781_25662# m1_20625_24224# m1_21729_25658# vss nfet$212
Xnfet$212_45 m1_15461_25858# m1_16085_25662# m1_15822_23922# vss nfet$212
Xnfet$212_34 m1_11278_25858# m1_13363_25658# m1_14156_24542# vss nfet$212
Xnfet$212_23 m1_11278_25858# vss m1_11415_25662# vss nfet$212
Xpfet$199_0 vdd m1_2590_19404# m1_2590_19404# m1_3458_19550# m1_n3534_17714# m1_n3534_17714#
+ pfet$199
Xnfet$215_9 sd5 vss m1_9331_15478# vss nfet$215
Xnfet$234_1 m1_n6433_17343# m1_n4377_15778# m1_n4994_16080# vss nfet$234
Xnfet$241_2 m1_n10933_25858# m1_n10309_25662# m1_n10572_23922# vss nfet$241
Xnfet$227_0 m1_31535_22102# m1_32818_21586# vss vss nfet$227
Xpfet$226_2 vdd m1_n5227_20152# vdd m1_n1927_20274# pfet$226
Xpfet$219_1 vdd vdd m1_n6111_25858# m1_n6856_24542# pfet$219
Xnfet$220_7 m1_25107_21786# vss m1_32193_25858# vss nfet$220
Xpfet$197_98 vdd m1_20104_16080# m1_19637_18030# m1_18665_17343# pfet$197
Xpfet$197_87 vdd vdd m1_18310_16080# m1_n7513_20152# pfet$197
Xpfet$197_76 vdd m1_17851_17714# vdd m1_18926_16202# pfet$197
Xpfet$197_65 vdd m1_24904_15778# m1_24287_16080# m1_23007_17836# pfet$197
Xpfet$197_21 vdd vdd m1_965_15478# sd7 pfet$197
Xpfet$197_10 vdd m1_8172_15778# m1_7555_16080# m1_6275_17836# pfet$197
Xpfet$197_32 vdd vdd m1_2905_18030# m1_3015_15778# pfet$197
Xpfet$197_43 vdd vdd m1_11271_18030# m1_11381_15778# pfet$197
Xpfet$197_54 vdd vdd m1_n1278_18030# m1_n1168_15778# pfet$197
Xnfet$213_6 m1_2384_21590# m1_2384_21590# m1_3871_22513# m1_3871_22513# m1_2843_21586#
+ vss nfet$213
Xpfet$205_7 vdd m1_32818_24542# vdd m1_33790_24346# pfet$205
Xnfet$220_12 m1_32675_25947# vss m1_28624_21786# vss nfet$220
Xpfet$197_109 vdd vdd m1_10299_17343# m1_13198_17714# pfet$197
Xnfet$211_3 m1_4509_24346# m1_4509_24346# m1_3394_25858# m1_3394_25858# m1_5456_25502#
+ vss nfet$211
Xnfet$215_78 m1_14641_17836# m1_15564_15778# m1_14743_16202# vss nfet$215
Xnfet$231_22 m1_15564_15778# m1_15564_15778# m1_15454_18030# m1_15454_18030# m1_15690_17358#
+ vss nfet$231
Xnfet$215_67 m1_17381_17714# vss m1_14482_17343# vss nfet$215
Xnfet$215_56 m1_24287_16080# vss m1_23930_15778# vss nfet$215
Xnfet$215_45 m1_n3064_17714# vss m1_n194_15778# vss nfet$215
Xnfet$215_34 m1_n2250_17343# vss m1_n2091_17836# vss nfet$215
Xnfet$215_23 m1_5302_17714# vss m1_4832_17714# vss nfet$215
Xnfet$215_12 m1_9485_17714# vss m1_12355_15778# vss nfet$215
Xnfet$231_11 m1_6377_16202# m1_6377_16202# vss vss m1_5859_16398# vss nfet$231
Xpfet$201_1 vdd vdd m1_n4377_15778# m1_n7247_17714# pfet$201
Xnfet$238_8 m1_9624_19404# m1_9624_19404# vss vss m1_n3724_21430# vss nfet$238
Xnfet$212_79 pd7 vss m1_19839_21786# vss nfet$212
Xnfet$212_68 m1_n7513_20152# vss m1_29607_24346# vss nfet$212
Xnfet$212_57 m1_20126_25858# vss m1_20268_25662# vss nfet$212
Xnfet$212_46 m1_20126_25858# vss m1_18073_21786# vss nfet$212
Xnfet$212_35 m1_15598_25662# m1_15822_23922# m1_16086_24542# vss nfet$212
Xnfet$212_24 m1_7095_25858# m1_7719_25662# m1_7456_23922# vss nfet$212
Xnfet$212_13 m1_11415_25662# m1_11639_23922# m1_11903_24542# vss nfet$212
Xpfet$199_1 vdd vdd vdd m1_2822_19850# m1_4620_20152# m1_4620_20152# pfet$199
Xnfet$234_2 m1_n6274_17836# m1_n5351_15778# m1_n6172_16202# vss nfet$234
Xpfet$226_3 vdd m1_n6839_20152# vdd m1_n927_19404# pfet$226
Xnfet$241_3 m1_n10796_25662# m1_n9952_24224# m1_n8848_25658# vss nfet$241
Xpfet$197_99 vdd m1_23109_16202# m1_22624_17518# m1_23007_17836# pfet$197
Xpfet$197_88 vdd vdd m1_18441_17518# m1_17851_17714# pfet$197
Xpfet$197_77 vdd vdd m1_17851_17714# m1_18310_16080# pfet$197
Xpfet$197_66 vdd vdd m1_24904_15778# m1_22034_17714# pfet$197
Xpfet$197_22 vdd vdd m1_3015_15778# m1_3372_16080# pfet$197
Xpfet$197_11 vdd vdd m1_9485_17714# m1_9944_16080# pfet$197
Xpfet$197_33 vdd vdd m1_5892_17518# m1_5302_17714# pfet$197
Xpfet$197_44 vdd vdd m1_649_17714# m1_1119_17714# pfet$197
Xpfet$197_55 vdd vdd m1_n2474_17518# m1_n3064_17714# pfet$197
Xnfet$220_8 m1_32193_25858# vss m1_32330_25662# vss nfet$220
Xnfet$213_7 m1_5771_21786# m1_5771_21786# m1_7388_22513# m1_7388_22513# m1_6992_21586#
+ vss nfet$213
Xnfet$220_13 m1_32675_25947# vss m1_32817_25662# vss nfet$220
Xpfet$224_0 vdd vdd vdd m1_n8047_19550# m1_n7513_20152# m1_n7513_20152# pfet$224
Xnfet$211_4 m1_12259_24224# m1_12259_24224# m1_11903_24542# m1_11903_24542# m1_12357_24542#
+ vss nfet$211
Xpfet$196_110 vdd m1_11903_24542# vdd m1_12875_24346# pfet$196
Xnfet$215_79 m1_15921_16080# vss m1_15564_15778# vss nfet$215
Xnfet$231_23 m1_18926_16202# m1_18926_16202# vss vss m1_18408_16398# vss nfet$231
Xnfet$215_68 m1_18665_17343# m1_18926_16202# m1_18441_17518# vss nfet$215
Xnfet$215_57 m1_22848_17343# m1_24904_15778# m1_24287_16080# vss nfet$215
Xnfet$215_46 m1_22034_17714# vss m1_21564_17714# vss nfet$215
Xnfet$215_24 m1_4832_17714# vss m1_1933_17343# vss nfet$215
Xnfet$215_13 m1_10458_17836# m1_11381_15778# m1_10560_16202# vss nfet$215
Xnfet$215_35 m1_n7513_20152# vss m1_5761_16080# vss nfet$215
Xnfet$231_12 m1_n1168_15778# m1_n1168_15778# m1_n1278_18030# m1_n1278_18030# m1_n1042_17358#
+ vss nfet$231
Xpfet$201_2 vdd vdd m1_n5351_15778# m1_n4994_16080# pfet$201
Xnfet$238_9 m1_n6380_21786# m1_n6380_21786# m1_n6839_21786# m1_n6839_21786# m1_n6282_21430#
+ vss nfet$238
Xnfet$212_69 m1_24309_25858# vss m1_26705_24542# vss nfet$212
Xnfet$212_58 m1_20005_23922# vss m1_20625_24224# vss nfet$212
Xnfet$212_47 m1_23964_25662# m1_24188_23922# m1_24452_24542# vss nfet$212
Xnfet$212_36 m1_11760_25858# vss m1_11039_21786# vss nfet$212
Xnfet$212_25 m1_7232_25662# m1_8076_24224# m1_9180_25658# vss nfet$212
Xnfet$212_14 m1_n7513_20152# vss m1_8692_24346# vss nfet$212
Xpfet$199_2 vdd m1_2590_19404# m1_2590_19404# m1_2822_19850# m1_2384_19550# m1_2384_19550#
+ pfet$199
Xnfet$234_3 m1_n6433_17343# m1_n6172_16202# m1_n6657_17518# vss nfet$234
Xnfet$241_4 m1_n4623_25487# m1_n2567_23922# m1_n3184_24224# vss nfet$241
Xpfet$197_89 vdd vdd m1_22848_17343# m1_25747_17714# pfet$197
Xpfet$197_78 vdd vdd m1_13514_15478# sd4 pfet$197
Xpfet$197_67 vdd m1_22034_17714# vdd m1_23109_16202# pfet$197
Xpfet$197_12 vdd m1_3989_15778# m1_3372_16080# m1_2092_17836# pfet$197
Xpfet$197_23 vdd m1_5302_17714# vdd m1_6377_16202# pfet$197
Xpfet$197_34 vdd vdd m1_5761_16080# m1_n7513_20152# pfet$197
Xpfet$197_45 vdd vdd m1_9944_16080# m1_n7513_20152# pfet$197
Xpfet$226_4 vdd vdd m1_n6839_20152# m1_n6973_21481# pfet$226
Xpfet$197_56 vdd m1_n1278_18030# vdd m1_n2605_16080# pfet$197
Xnfet$220_9 m1_n7513_20152# vss m1_33790_24346# vss nfet$220
Xnfet$213_8 m1_23486_21590# m1_23486_21590# m1_24973_22513# m1_24973_22513# m1_23945_21586#
+ vss nfet$213
Xnfet$232_0 m1_4620_20152# m1_4620_20152# m1_2590_19404# m1_2590_19404# m1_3454_20470#
+ vss nfet$232
Xpfet$224_1 vdd m1_n8283_19850# m1_n8283_19850# m1_n8047_19550# m1_n8283_20611# m1_n8283_20611#
+ pfet$224
Xpfet$217_0 vdd vdd vdd m1_n6624_23622# m1_n7082_23622# m1_n7082_23622# pfet$217
Xnfet$211_5 m1_8692_24346# m1_8692_24346# vss vss m1_8174_24542# vss nfet$211
Xpfet$196_100 vdd vdd m1_29607_24346# m1_n7513_20152# pfet$196
Xnfet$215_58 m1_23007_17836# m1_23930_15778# m1_23109_16202# vss nfet$215
Xnfet$215_47 m1_22034_17714# vss m1_22624_17518# vss nfet$215
Xnfet$215_25 m1_2092_17836# m1_3372_16080# m1_2905_18030# vss nfet$215
Xnfet$215_14 m1_6116_17343# m1_8172_15778# m1_7555_16080# vss nfet$215
Xnfet$215_36 m1_n3064_17714# vss m1_n2474_17518# vss nfet$215
Xnfet$231_24 m1_18310_16080# m1_18310_16080# m1_17851_17714# m1_17851_17714# m1_18408_16398#
+ vss nfet$231
Xnfet$215_69 m1_17851_17714# vss m1_17381_17714# vss nfet$215
Xnfet$231_13 m1_n2605_16080# m1_n2605_16080# vss vss m1_n1042_17358# vss nfet$231
Xpfet$201_3 vdd vdd m1_n6657_17518# m1_n7247_17714# pfet$201
Xnfet$212_59 m1_19644_25858# m1_20268_25662# m1_20005_23922# vss nfet$212
Xnfet$212_48 m1_18073_21786# vss m1_23827_25858# vss nfet$212
Xnfet$212_37 m1_11039_21786# vss m1_15461_25858# vss nfet$212
Xnfet$212_26 m1_7095_25858# m1_9180_25658# m1_9973_24542# vss nfet$212
Xnfet$212_15 m1_7232_25662# m1_7456_23922# m1_7720_24542# vss nfet$212
Xpfet$200_10 vdd vdd m1_23486_21590# m1_23356_21786# pfet$200
Xpfet$199_3 vdd vdd vdd m1_3458_19550# m1_n3218_15478# m1_n3218_15478# pfet$199
Xnfet$234_4 m1_27031_17343# m1_27292_16202# m1_26807_17518# vss nfet$234
Xnfet$241_5 m1_n4464_25980# m1_n3541_23922# m1_n4362_24346# vss nfet$241
Xpfet$197_79 vdd m1_15564_15778# m1_14743_16202# m1_14482_17343# pfet$197
Xpfet$197_68 vdd vdd m1_22034_17714# m1_22493_16080# pfet$197
Xpfet$197_13 vdd vdd m1_5148_15478# sd6 pfet$197
Xpfet$197_0 vdd vdd m1_12355_15778# m1_9485_17714# pfet$197
Xpfet$197_24 vdd m1_6377_16202# m1_5892_17518# m1_6275_17836# pfet$197
Xpfet$197_35 vdd vdd m1_9015_17714# m1_9485_17714# pfet$197
Xpfet$197_46 vdd vdd m1_n2250_17343# m1_649_17714# pfet$197
Xpfet$197_57 vdd m1_n1989_16202# m1_n2474_17518# m1_n2091_17836# pfet$197
Xnfet$213_9 m1_23356_21786# m1_23356_21786# m1_24973_22513# m1_24973_22513# m1_24577_21586#
+ vss nfet$213
Xnfet$225_0 m1_21456_22513# m1_21456_22513# m1_30256_19792# m1_30256_19792# m1_30492_20470#
+ vss nfet$225
Xnfet$232_1 m1_1103_20152# m1_1103_20152# m1_n927_19404# m1_n927_19404# m1_n63_20470#
+ vss nfet$232
Xpfet$224_2 vdd m1_n8283_20611# m1_n8283_20611# m1_n8047_22344# m1_n8145_21908# m1_n8145_21908#
+ pfet$224
Xpfet$217_1 vdd m1_n6856_24542# m1_n6856_24542# m1_n6624_23622# m1_n8283_19850# m1_n8283_19850#
+ pfet$217
Xpfet$196_101 vdd vdd m1_28010_25858# m1_21590_21786# pfet$196
Xnfet$211_6 m1_8076_24224# m1_8076_24224# m1_7720_24542# m1_7720_24542# m1_8174_24542#
+ vss nfet$211
Xnfet$231_25 m1_14743_16202# m1_14743_16202# vss vss m1_14225_16398# vss nfet$231
Xnfet$215_59 m1_17851_17714# vss m1_20721_15778# vss nfet$215
Xnfet$215_48 m1_18824_17836# m1_20104_16080# m1_19637_18030# vss nfet$215
Xnfet$215_26 m1_5302_17714# vss m1_5892_17518# vss nfet$215
Xnfet$215_15 m1_5302_17714# vss m1_8172_15778# vss nfet$215
Xnfet$215_37 m1_n7513_20152# vss m1_n2605_16080# vss nfet$215
Xnfet$231_14 m1_n2605_16080# m1_n2605_16080# m1_n3064_17714# m1_n3064_17714# m1_n2507_16398#
+ vss nfet$231
Xpfet$201_4 vdd vdd m1_n6433_17343# m1_n3534_17714# pfet$201
Xnfet$212_49 m1_19781_25662# m1_20005_23922# m1_20269_24542# vss nfet$212
Xnfet$212_38 m1_n7513_20152# vss m1_12875_24346# vss nfet$212
Xnfet$212_27 m1_7577_25858# vss m1_7719_25662# vss nfet$212
Xnfet$212_16 m1_4005_21786# vss m1_7095_25858# vss nfet$212
Xpfet$200_11 vdd vdd m1_18705_21786# m1_18073_21786# pfet$200
Xpfet$199_4 vdd m1_6107_19404# m1_6107_19404# m1_6339_19850# m1_5901_19550# m1_5901_19550#
+ pfet$199
Xnfet$234_5 m1_27031_17343# m1_29087_15778# m1_28470_16080# vss nfet$234
Xnfet$241_6 m1_n4464_25980# m1_n3184_24224# m1_n3651_26174# vss nfet$241
Xpfet$197_14 vdd vdd m1_2092_17836# m1_1933_17343# pfet$197
Xpfet$197_1 vdd vdd m1_11381_15778# m1_11738_16080# pfet$197
Xpfet$197_25 vdd vdd m1_1709_17518# m1_1119_17714# pfet$197
Xpfet$197_36 vdd vdd m1_6116_17343# m1_9015_17714# pfet$197
Xpfet$197_69 vdd vdd m1_20721_15778# m1_17851_17714# pfet$197
Xpfet$197_47 vdd m1_11738_16080# m1_11271_18030# m1_10299_17343# pfet$197
Xpfet$197_58 vdd vdd m1_n3534_17714# m1_n3064_17714# pfet$197
Xnfet$225_1 m1_14422_22513# m1_14422_22513# m1_31535_19792# m1_31535_19792# m1_31771_20470#
+ vss nfet$225
Xnfet$232_2 m1_n3218_15478# m1_n3218_15478# m1_2590_19404# m1_2590_19404# m1_2822_20470#
+ vss nfet$232
Xnfet$218_0 sd9 vss m1_n7401_15478# vss nfet$218
Xpfet$224_3 vdd vdd vdd m1_n8047_22344# m1_n8283_19850# m1_n8283_19850# pfet$224
Xnfet$211_7 m1_9180_25658# m1_9180_25658# vss vss m1_9639_25502# vss nfet$211
Xpfet$196_102 vdd m1_28371_23922# m1_28635_24542# m1_28010_25858# pfet$196
Xnfet$231_26 m1_14127_16080# m1_14127_16080# m1_13668_17714# m1_13668_17714# m1_14225_16398#
+ vss nfet$231
Xnfet$215_49 m1_21564_17714# vss m1_18665_17343# vss nfet$215
Xnfet$215_27 m1_1119_17714# vss m1_3989_15778# vss nfet$215
Xnfet$215_16 m1_6275_17836# m1_7198_15778# m1_6377_16202# vss nfet$215
Xnfet$215_38 m1_n2250_17343# m1_n1989_16202# m1_n2474_17518# vss nfet$215
Xnfet$231_15 m1_n1989_16202# m1_n1989_16202# vss vss m1_n2507_16398# vss nfet$231
Xpfet$222_0 vdd vdd m1_n10796_25662# m1_n10933_25858# pfet$222
Xpfet$201_5 vdd vdd m1_n6788_16080# m1_n7513_20152# pfet$201
Xnfet$212_28 m1_3394_25858# vss m1_4005_21786# vss nfet$212
Xnfet$212_17 m1_11639_23922# vss m1_12259_24224# vss nfet$212
Xnfet$212_39 pd4 vss m1_9288_21786# vss nfet$212
Xpfet$200_12 vdd vdd m1_16452_21590# m1_16322_21786# pfet$200
Xpfet$199_5 vdd vdd vdd m1_n695_19850# m1_1103_20152# m1_1103_20152# pfet$199
Xnfet$234_6 m1_27190_17836# m1_28113_15778# m1_27292_16202# vss nfet$234
Xnfet$241_7 m1_n4623_25487# m1_n4362_24346# m1_n4847_25662# vss nfet$241
Xpfet$197_15 vdd vdd m1_5302_17714# m1_5761_16080# pfet$197
Xpfet$197_2 vdd m1_12355_15778# m1_11738_16080# m1_10458_17836# pfet$197
Xpfet$197_26 vdd vdd m1_4832_17714# m1_5302_17714# pfet$197
Xpfet$197_37 vdd m1_7555_16080# m1_7088_18030# m1_6116_17343# pfet$197
Xpfet$197_48 vdd vdd m1_n3064_17714# m1_n2605_16080# pfet$197
Xpfet$197_59 vdd vdd m1_n2605_16080# m1_n7513_20152# pfet$197
Xnfet$218_1 sd2 vss m1_21880_15478# vss nfet$218
Xnfet$225_2 m1_17939_22513# m1_17939_22513# vss vss m1_31771_20470# vss nfet$225
Xnfet$232_3 m1_8137_20152# m1_8137_20152# m1_6107_19404# m1_6107_19404# m1_6971_20470#
+ vss nfet$232
Xpfet$222_10 vdd vdd m1_n10933_25858# fin pfet$222
Xnfet$211_8 m1_8692_24346# m1_8692_24346# m1_7577_25858# m1_7577_25858# m1_9639_25502#
+ vss nfet$211
Xpfet$196_103 vdd vdd m1_28635_24542# m1_28991_24224# pfet$196
Xnfet$230_0 fout vss m1_35837_22102# vss nfet$230
Xnfet$231_27 m1_18310_16080# m1_18310_16080# vss vss m1_19873_17358# vss nfet$231
Xnfet$231_16 m1_19747_15778# m1_19747_15778# m1_19637_18030# m1_19637_18030# m1_19873_17358#
+ vss nfet$231
Xnfet$215_28 m1_1933_17343# vss m1_2092_17836# vss nfet$215
Xnfet$215_17 m1_649_17714# vss m1_n2250_17343# vss nfet$215
Xnfet$215_39 m1_n3064_17714# vss m1_n3534_17714# vss nfet$215
Xpfet$222_1 vdd vdd m1_n10309_25662# m1_n10452_25858# pfet$222
Xpfet$215_0 vdd m1_n4377_15778# m1_n4994_16080# m1_n6274_17836# pfet$215
Xpfet$201_6 vdd vdd m1_n7383_17599# m1_n7247_17714# pfet$201
Xnfet$212_29 m1_15943_25858# vss m1_14556_21786# vss nfet$212
Xnfet$212_18 m1_7095_25858# vss m1_7232_25662# vss nfet$212
Xpfet$200_13 vdd vdd m1_15188_21786# m1_14556_21786# pfet$200
Xpfet$199_6 vdd vdd vdd m1_6339_19850# m1_8137_20152# m1_8137_20152# pfet$199
Xnfet$234_7 m1_27190_17836# m1_28470_16080# m1_28003_18030# vss nfet$234
Xpfet$197_16 vdd vdd m1_3989_15778# m1_1119_17714# pfet$197
Xpfet$197_3 vdd m1_11381_15778# m1_10560_16202# m1_10299_17343# pfet$197
Xpfet$197_27 vdd m1_2194_16202# m1_1709_17518# m1_2092_17836# pfet$197
Xpfet$197_38 vdd vdd m1_7088_18030# m1_7198_15778# pfet$197
Xpfet$197_49 vdd m1_n194_15778# m1_n811_16080# m1_n2091_17836# pfet$197
Xnfet$218_2 sd1 vss m1_26063_15478# vss nfet$218
Xnfet$225_3 m1_24973_22513# m1_24973_22513# vss vss m1_30492_20470# vss nfet$225
Xnfet$232_4 m1_965_15478# m1_965_15478# m1_6107_19404# m1_6107_19404# m1_6339_20470#
+ vss nfet$232
Xpfet$222_11 vdd vdd m1_n9336_24346# vss pfet$222
Xnfet$211_9 m1_17058_24346# m1_17058_24346# vss vss m1_16540_24542# vss nfet$211
Xpfet$196_104 vdd m1_25912_25658# m1_26705_24542# m1_23964_25662# pfet$196
Xnfet$230_1 define m1_35837_22102# vss vss nfet$230
Xnfet$231_17 m1_22493_16080# m1_22493_16080# vss vss m1_24056_17358# vss nfet$231
Xnfet$215_29 m1_3372_16080# vss m1_3015_15778# vss nfet$215
Xnfet$215_18 m1_1119_17714# vss m1_649_17714# vss nfet$215
Xnfet$223_0 m1_n290_24224# m1_n290_24224# m1_n646_24542# m1_n646_24542# m1_n192_24542#
+ vss nfet$223
Xpfet$215_1 vdd m1_n5351_15778# m1_n6172_16202# m1_n6433_17343# pfet$215
Xpfet$222_2 vdd vdd m1_n9952_24224# m1_n10572_23922# pfet$222
Xpfet$208_0 vdd m1_n647_25662# m1_n910_23922# m1_n1134_25662# pfet$208
Xpfet$201_7 vdd vdd m1_27190_17836# m1_27031_17343# pfet$201
Xnfet$212_19 m1_7456_23922# vss m1_8076_24224# vss nfet$212
Xpfet$200_14 vdd vdd m1_19969_21590# m1_19839_21786# pfet$200
Xpfet$199_7 vdd vdd vdd m1_6975_19550# m1_965_15478# m1_965_15478# pfet$199
Xpfet$197_17 vdd vdd m1_n2091_17836# m1_n2250_17343# pfet$197
Xpfet$197_4 vdd m1_9485_17714# vdd m1_10560_16202# pfet$197
Xpfet$197_28 vdd m1_2905_18030# vdd m1_1578_16080# pfet$197
Xpfet$197_39 vdd m1_7088_18030# vdd m1_5761_16080# pfet$197
Xnfet$225_4 m1_32818_20470# m1_32818_20470# vss vss m1_34329_20470# vss nfet$225
Xnfet$232_5 m1_5148_15478# m1_5148_15478# m1_9624_19404# m1_9624_19404# m1_9856_20470#
+ vss nfet$232
Xpfet$222_12 vdd vdd m1_n7082_23622# m1_n8625_26174# pfet$222
Xpfet$196_105 vdd vdd m1_30888_24542# m1_28492_25858# pfet$196
Xnfet$223_1 m1_814_25658# m1_814_25658# vss vss m1_1273_25502# vss nfet$223
Xnfet$215_19 m1_n7513_20152# vss m1_1578_16080# vss nfet$215
Xnfet$216_0 m1_n1263_21786# vss m1_n1133_21590# vss nfet$216
Xnfet$231_18 m1_23930_15778# m1_23930_15778# m1_23820_18030# m1_23820_18030# m1_24056_17358#
+ vss nfet$231
Xpfet$215_2 vdd m1_n4994_16080# m1_n5461_18030# m1_n6433_17343# pfet$215
Xpfet$222_3 vdd vdd m1_n4978_24224# vss pfet$222
Xpfet$208_1 vdd m1_n910_23922# m1_n646_24542# m1_n1271_25858# pfet$208
Xpfet$201_8 vdd vdd m1_28113_15778# m1_28470_16080# pfet$201
Xpfet$220_0 vdd vdd m1_n8625_26174# m1_n9336_24346# pfet$220
Xpfet$200_15 vdd vdd m1_27003_21590# m1_26873_21786# pfet$200
Xpfet$199_8 vdd m1_9624_19404# m1_9624_19404# m1_10492_19550# m1_4832_17714# m1_4832_17714#
+ pfet$199
Xpfet$197_18 vdd m1_1119_17714# vdd m1_2194_16202# pfet$197
Xpfet$197_5 vdd m1_7198_15778# m1_6377_16202# m1_6116_17343# pfet$197
Xpfet$197_29 vdd vdd m1_1578_16080# m1_n7513_20152# pfet$197
Xnfet$246_0 m1_n4485_20152# m1_n6380_21786# vss vss nfet$246
Xnfet$225_5 m1_32818_21586# m1_32818_21586# m1_34093_19792# m1_34093_19792# m1_34329_20470#
+ vss nfet$225
Xnfet$232_6 m1_11654_20152# m1_11654_20152# m1_9624_19404# m1_9624_19404# m1_10488_20470#
+ vss nfet$232
Xpfet$222_13 vdd vdd m1_n8055_24542# m1_n8625_26174# pfet$222
Xpfet$196_106 vdd vdd m1_25107_21786# m1_28492_25858# pfet$196
Xnfet$223_2 m1_326_24346# m1_326_24346# m1_n789_25858# m1_n789_25858# m1_1273_25502#
+ vss nfet$223
Xnfet$231_19 m1_23109_16202# m1_23109_16202# vss vss m1_22591_16398# vss nfet$231
Xpfet$215_3 vdd m1_n6172_16202# m1_n6657_17518# m1_n6274_17836# pfet$215
Xpfet$222_4 vdd vdd m1_n5571_25662# m1_n10452_25858# pfet$222
Xnfet$216_1 m1_11039_21786# vss m1_11671_21786# vss nfet$216
Xpfet$208_2 vdd m1_n290_24224# m1_814_25658# m1_n1271_25858# pfet$208
Xpfet$201_9 vdd vdd m1_29087_15778# m1_26217_17714# pfet$201
Xpfet$213_0 vdd m1_32818_20470# m1_32818_20470# m1_33050_19550# m1_30256_19792# m1_30256_19792#
+ pfet$213
Xpfet$220_1 vdd m1_n8625_26174# vdd m1_n8848_25658# pfet$220
Xpfet$200_16 vdd vdd m1_29256_21786# m1_28624_21786# pfet$200
Xpfet$199_9 vdd m1_9624_19404# m1_9624_19404# m1_9856_19850# m1_9418_19550# m1_9418_19550#
+ pfet$199
Xpfet$197_19 vdd m1_3015_15778# m1_2194_16202# m1_1933_17343# pfet$197
Xpfet$197_6 vdd vdd m1_7198_15778# m1_7555_16080# pfet$197
Xnfet$246_1 m1_n5227_20152# vss m1_n6380_21786# vss nfet$246
Xnfet$239_0 m1_n8625_26174# vss m1_n8055_24542# vss nfet$239
Xnfet$225_6 m1_354_22513# m1_354_22513# m1_31535_22102# m1_31535_22102# m1_31771_21430#
+ vss nfet$225
Xnfet$232_7 m1_n7401_15478# m1_n7401_15478# m1_n927_19404# m1_n927_19404# m1_n695_20470#
+ vss nfet$232
Xpfet$196_107 vdd m1_24309_25858# vdd m1_25912_25658# pfet$196
Xpfet$215_4 vdd m1_28113_15778# m1_27292_16202# m1_27031_17343# pfet$215
Xnfet$223_3 m1_326_24346# m1_326_24346# vss vss m1_n192_24542# vss nfet$223
Xpfet$208_3 vdd m1_814_25658# m1_1607_24542# m1_n1134_25662# pfet$208
Xpfet$222_5 vdd vdd m1_n4847_25662# m1_n10452_25858# pfet$222
Xnfet$216_2 m1_12805_21786# vss m1_12935_21590# vss nfet$216
Xnfet$221_0 m1_n1134_25662# m1_n910_23922# m1_n646_24542# vss nfet$221
Xpfet$206_0 vdd vdd vdd m1_33050_22344# m1_31535_22102# m1_31535_22102# pfet$206
Xpfet$213_1 vdd vdd vdd m1_33050_19550# m1_31535_19792# m1_31535_19792# pfet$213
Xpfet$220_2 vdd m1_n3651_26174# vdd m1_n4978_24224# pfet$220
Xpfet$200_17 vdd vdd m1_25739_21786# m1_25107_21786# pfet$200
Xnfet$213_10 m1_19839_21786# m1_19839_21786# m1_21456_22513# m1_21456_22513# m1_21060_21586#
+ vss nfet$213
Xnfet$239_1 m1_n8625_26174# vss m1_n7082_23622# vss nfet$239
Xpfet$197_7 vdd vdd m1_6275_17836# m1_6116_17343# pfet$197
Xnfet$225_7 m1_3871_22513# m1_3871_22513# vss vss m1_31771_21430# vss nfet$225
Xnfet$232_8 m1_26063_15478# m1_26063_15478# m1_n3822_20130# m1_n3822_20130# m1_27441_20470#
+ vss nfet$232
Xpfet$198_30 vdd vdd vdd m1_17539_22402# m1_16322_21786# m1_16322_21786# pfet$198
Xpfet$196_108 vdd vdd m1_25424_24346# m1_n7513_20152# pfet$196
Xnfet$223_4 m1_33174_24224# m1_33174_24224# m1_32818_24542# m1_32818_24542# m1_33272_24542#
+ vss nfet$223
Xpfet$222_6 vdd vdd m1_n4623_25487# fin pfet$222
Xnfet$216_3 m1_9288_21786# vss m1_9418_21590# vss nfet$216
Xpfet$208_4 vdd m1_33174_24224# m1_34278_25658# m1_32193_25858# pfet$208
Xpfet$215_5 vdd m1_29087_15778# m1_28470_16080# m1_27190_17836# pfet$215
Xpfet$213_2 vdd m1_32818_21586# m1_32818_21586# m1_33050_22344# m1_30256_22102# m1_30256_22102#
+ pfet$213
Xnfet$216_10 m1_21590_21786# vss m1_22222_21786# vss nfet$216
Xnfet$214_0 m1_n3534_17714# m1_n3534_17714# vss vss m1_3454_20470# vss nfet$214
Xnfet$221_1 m1_n1271_25858# m1_n647_25662# m1_n910_23922# vss nfet$221
Xpfet$220_3 vdd vdd m1_n3651_26174# m1_n3541_23922# pfet$220
Xnfet$213_11 m1_19969_21590# m1_19969_21590# m1_21456_22513# m1_21456_22513# m1_20428_21586#
+ vss nfet$213
Xpfet$197_8 vdd vdd m1_9331_15478# sd5 pfet$197
Xnfet$239_2 vss vss m1_n9336_24346# vss nfet$239
Xnfet$224_10 m1_21590_21786# m1_21590_21786# vss vss m1_20428_21586# vss nfet$224
Xnfet$232_9 m1_29239_20152# m1_29239_20152# m1_n3822_20130# m1_n3822_20130# m1_28073_20470#
+ vss nfet$232
Xnfet$244_0 m1_n4485_21904# m1_n5764_21786# vss vss nfet$244
Xpfet$198_31 vdd vdd vdd m1_27462_22102# m1_27003_21590# m1_27003_21590# pfet$198
Xpfet$198_20 vdd vdd vdd m1_20428_22102# m1_19969_21590# m1_19969_21590# pfet$198
Xnfet$219_10 m1_26217_17714# vss m1_29087_15778# vss nfet$219
Xpfet$196_109 vdd m1_12259_24224# m1_13363_25658# m1_11278_25858# pfet$196
Xnfet$223_5 m1_33790_24346# m1_33790_24346# vss vss m1_33272_24542# vss nfet$223
Xnfet$216_4 m1_7522_21786# vss m1_8154_21786# vss nfet$216
Xpfet$208_5 vdd m1_32817_25662# m1_32554_23922# m1_32330_25662# pfet$208
Xpfet$215_6 vdd m1_28470_16080# m1_28003_18030# m1_27031_17343# pfet$215
Xpfet$222_7 vdd vdd m1_n3541_23922# m1_n3184_24224# pfet$222
Xnfet$214_1 m1_2384_19550# m1_2384_19550# vss vss m1_2822_20470# vss nfet$214
Xpfet$220_4 vdd m1_n10452_25858# vdd m1_n4362_24346# pfet$220
Xnfet$221_2 m1_n1271_25858# m1_814_25658# m1_1607_24542# vss nfet$221
Xnfet$216_11 m1_18073_21786# vss m1_18705_21786# vss nfet$216
Xnfet$232_10 m1_9331_15478# m1_9331_15478# m1_n3822_21786# m1_n3822_21786# m1_13373_20470#
+ vss nfet$232
Xpfet$211_0 vdd vdd vdd m1_36073_22344# define define pfet$211
Xnfet$213_12 m1_16322_21786# m1_16322_21786# m1_17939_22513# m1_17939_22513# m1_17543_21586#
+ vss nfet$213
Xpfet$197_9 vdd vdd m1_8172_15778# m1_5302_17714# pfet$197
Xnfet$239_3 fin vss m1_n10933_25858# vss nfet$239
Xnfet$224_11 m1_22222_21786# m1_22222_21786# vss vss m1_21060_21586# vss nfet$224
Xnfet$244_1 m1_n5227_21418# vss m1_n5764_21786# vss nfet$244
Xnfet$237_0 m1_n7082_23622# m1_n6856_24542# vss vss nfet$237
Xnfet$219_11 m1_27031_17343# vss m1_27190_17836# vss nfet$219
Xnfet$223_6 m1_33790_24346# m1_33790_24346# m1_32675_25947# m1_32675_25947# m1_34737_25502#
+ vss nfet$223
Xpfet$198_32 vdd m1_28490_22513# m1_28490_22513# m1_28090_22402# m1_28624_21786# m1_28624_21786#
+ pfet$198
Xpfet$198_21 vdd vdd vdd m1_21056_22402# m1_19839_21786# m1_19839_21786# pfet$198
Xnfet$216_5 m1_488_21786# vss m1_1120_21786# vss nfet$216
Xpfet$198_10 vdd m1_3871_22513# m1_3871_22513# m1_2843_22102# m1_4637_21786# m1_4637_21786#
+ pfet$198
Xpfet$208_6 vdd m1_34278_25658# m1_35071_24542# m1_32330_25662# pfet$208
Xpfet$215_7 vdd m1_27292_16202# m1_26807_17518# m1_27190_17836# pfet$215
Xpfet$222_8 vdd vdd m1_n2567_23922# m1_n7320_25516# pfet$222
Xnfet$221_3 m1_n1134_25662# m1_n290_24224# m1_814_25658# vss nfet$221
Xnfet$214_2 m1_5901_19550# m1_5901_19550# vss vss m1_6339_20470# vss nfet$214
Xnfet$216_12 m1_14556_21786# vss m1_15188_21786# vss nfet$216
Xnfet$232_11 m1_15171_20152# m1_15171_20152# m1_n3822_21786# m1_n3822_21786# m1_14005_20470#
+ vss nfet$232
Xpfet$220_5 vdd vdd m1_n10308_24542# m1_n9952_24224# pfet$220
Xpfet$211_1 vdd m1_35837_22102# m1_35837_22102# m1_36073_22344# fout fout pfet$211
Xpfet$204_0 vdd vdd m1_n647_25662# m1_n789_25858# pfet$204
Xnfet$213_13 m1_16452_21590# m1_16452_21590# m1_17939_22513# m1_17939_22513# m1_16911_21586#
+ vss nfet$213
Xnfet$239_4 m1_n10572_23922# vss m1_n9952_24224# vss nfet$239
Xnfet$224_12 m1_18073_21786# m1_18073_21786# vss vss m1_16911_21586# vss nfet$224
Xnfet$219_12 m1_28470_16080# vss m1_28113_15778# vss nfet$219
Xnfet$244_2 m1_n6839_21786# vss m1_n6973_21481# vss nfet$244
Xnfet$237_1 m1_n8283_19850# vss m1_n6856_24542# vss nfet$237
Xnfet$223_7 m1_34278_25658# m1_34278_25658# vss vss m1_34737_25502# vss nfet$223
Xpfet$198_33 vdd m1_28490_22513# m1_28490_22513# m1_27462_22102# m1_29256_21786# m1_29256_21786#
+ pfet$198
Xpfet$198_22 vdd m1_21456_22513# m1_21456_22513# m1_20428_22102# m1_22222_21786# m1_22222_21786#
+ pfet$198
Xpfet$198_11 vdd vdd vdd m1_2843_22102# m1_2384_21590# m1_2384_21590# pfet$198
Xpfet$208_7 vdd m1_32554_23922# m1_32818_24542# m1_32193_25858# pfet$208
Xpfet$222_9 vdd vdd m1_n4464_25980# m1_n4623_25487# pfet$222
Xnfet$216_6 m1_5771_21786# vss m1_5901_21590# vss nfet$216
Xnfet$221_4 m1_32193_25858# m1_34278_25658# m1_35071_24542# vss nfet$221
Xnfet$214_3 m1_4832_17714# m1_4832_17714# vss vss m1_10488_20470# vss nfet$214
Xnfet$216_13 m1_16322_21786# vss m1_16452_21590# vss nfet$216
Xnfet$232_12 m1_18688_20152# m1_18688_20152# m1_n1927_20274# m1_n1927_20274# m1_17522_20470#
+ vss nfet$232
Xpfet$220_6 vdd m1_n10308_24542# vdd m1_n9336_24346# pfet$220
Xnfet$212_0 m1_3394_25858# vss m1_5790_24542# vss nfet$212
Xpfet$204_1 vdd vdd m1_n1134_25662# m1_n1271_25858# pfet$204
Xnfet$213_14 m1_12805_21786# m1_12805_21786# m1_14422_22513# m1_14422_22513# m1_14026_21586#
+ vss nfet$213
Xnfet$239_5 m1_n10933_25858# vss m1_n10796_25662# vss nfet$239
Xnfet$224_13 m1_18705_21786# m1_18705_21786# vss vss m1_17543_21586# vss nfet$224
Xnfet$219_13 m1_26217_17714# vss m1_25747_17714# vss nfet$219
Xpfet$198_34 vdd vdd vdd m1_28090_22402# m1_26873_21786# m1_26873_21786# pfet$198
Xpfet$198_23 vdd vdd vdd m1_23945_22102# m1_23486_21590# m1_23486_21590# pfet$198
Xpfet$198_12 vdd vdd vdd m1_3471_22402# m1_2254_21786# m1_2254_21786# pfet$198
Xnfet$242_0 m1_n7186_25858# vss m1_n7320_25516# vss nfet$242
Xnfet$216_7 m1_4005_21786# vss m1_4637_21786# vss nfet$216
Xpfet$227_0 vdd vdd vdd m1_n5019_19550# m1_n4485_20152# m1_n4485_20152# pfet$227
Xnfet$221_5 m1_32330_25662# m1_33174_24224# m1_34278_25658# vss nfet$221
Xnfet$214_4 m1_9418_19550# m1_9418_19550# vss vss m1_9856_20470# vss nfet$214
Xnfet$216_14 m1_19839_21786# vss m1_19969_21590# vss nfet$216
Xnfet$232_13 m1_13514_15478# m1_13514_15478# m1_n1927_20274# m1_n1927_20274# m1_16890_20470#
+ vss nfet$232
Xpfet$220_7 vdd vdd m1_n10452_25858# m1_n4978_24224# pfet$220
Xnfet$212_1 m1_2912_25858# m1_4997_25658# m1_5790_24542# vss nfet$212
Xpfet$204_2 vdd vdd m1_n1271_25858# m1_n10452_25858# pfet$204
Xnfet$213_15 m1_26873_21786# m1_26873_21786# m1_28490_22513# m1_28490_22513# m1_28094_21586#
+ vss nfet$213
Xnfet$239_6 m1_n10452_25858# vss m1_n10309_25662# vss nfet$239
Xnfet$224_14 m1_15188_21786# m1_15188_21786# vss vss m1_14026_21586# vss nfet$224
Xpfet$201_10 vdd vdd m1_27031_17343# m1_n10452_25858# pfet$201
Xpfet$198_35 vdd vdd vdd m1_13394_22102# m1_12935_21590# m1_12935_21590# pfet$198
Xpfet$198_24 vdd m1_17939_22513# m1_17939_22513# m1_16911_22102# m1_18705_21786# m1_18705_21786#
+ pfet$198
Xpfet$198_13 vdd vdd vdd m1_6988_22402# m1_5771_21786# m1_5771_21786# pfet$198
Xnfet$216_8 m1_2254_21786# vss m1_2384_21590# vss nfet$216
Xnfet$235_0 m1_n5351_15778# m1_n5351_15778# m1_n5461_18030# m1_n5461_18030# m1_n5225_17358#
+ vss nfet$235
Xnfet$242_1 m1_n6856_24542# vss m1_n6111_25858# vss nfet$242
Xnfet$221_6 m1_32193_25858# m1_32817_25662# m1_32554_23922# vss nfet$221
Xnfet$216_15 m1_28624_21786# vss m1_29256_21786# vss nfet$216
Xnfet$214_5 m1_649_17714# m1_649_17714# vss vss m1_6971_20470# vss nfet$214
Xnfet$232_14 m1_22205_20152# m1_22205_20152# m1_n2543_20130# m1_n2543_20130# m1_21039_20470#
+ vss nfet$232
Xpfet$204_10 vdd vdd m1_35071_24542# m1_32675_25947# pfet$204
Xnfet$212_2 m1_n7513_20152# vss m1_4509_24346# vss nfet$212
Xpfet$204_3 vdd vdd m1_1607_24542# m1_n789_25858# pfet$204
Xpfet$196_90 vdd vdd m1_24309_25858# m1_25424_24346# pfet$196
Xnfet$213_16 m1_27003_21590# m1_27003_21590# m1_28490_22513# m1_28490_22513# m1_27462_21586#
+ vss nfet$213
Xpfet$202_0 vdd vdd m1_2384_19550# m1_n3534_17714# pfet$202
Xpfet$201_11 vdd vdd m1_26807_17518# m1_26217_17714# pfet$201
Xnfet$239_7 m1_n7320_25516# vss m1_n2567_23922# vss nfet$239
Xnfet$224_15 m1_14556_21786# m1_14556_21786# vss vss m1_13394_21586# vss nfet$224
Xpfet$198_25 vdd m1_17939_22513# m1_17939_22513# m1_17539_22402# m1_18073_21786# m1_18073_21786#
+ pfet$198
Xpfet$198_14 vdd vdd vdd m1_n46_22402# m1_n1263_21786# m1_n1263_21786# pfet$198
Xnfet$216_9 m1_23356_21786# vss m1_23486_21590# vss nfet$216
Xnfet$228_0 m1_34093_19792# vss m1_34843_21786# vss nfet$228
Xnfet$235_1 m1_n6788_16080# m1_n6788_16080# vss vss m1_n5225_17358# vss nfet$235
Xnfet$221_7 m1_32330_25662# m1_32554_23922# m1_32818_24542# vss nfet$221
Xnfet$214_6 m1_n1133_19550# m1_n1133_19550# vss vss m1_n695_20470# vss nfet$214
Xnfet$216_16 m1_26873_21786# vss m1_27003_21590# vss nfet$216
Xnfet$232_15 m1_17697_15478# m1_17697_15478# m1_n2543_20130# m1_n2543_20130# m1_20407_20470#
+ vss nfet$232
Xpfet$204_11 vdd vdd m1_32817_25662# m1_32675_25947# pfet$204
Xnfet$212_3 m1_488_21786# vss m1_2912_25858# vss nfet$212
Xpfet$204_4 vdd vdd m1_488_21786# m1_n789_25858# pfet$204
Xnfet$213_17 m1_12935_21590# m1_12935_21590# m1_14422_22513# m1_14422_22513# m1_13394_21586#
+ vss nfet$213
Xpfet$196_91 vdd vdd m1_23356_21786# pd8 pfet$196
Xpfet$196_80 vdd vdd m1_17058_24346# m1_n7513_20152# pfet$196
Xpfet$202_1 vdd vdd m1_4620_20152# m1_n3218_15478# pfet$202
Xpfet$201_12 vdd vdd m1_26676_16080# m1_n7513_20152# pfet$201
Xnfet$239_8 m1_n4623_25487# vss m1_n4464_25980# vss nfet$239
Xnfet$224_16 m1_28624_21786# m1_28624_21786# vss vss m1_27462_21586# vss nfet$224
Xpfet$198_26 vdd vdd vdd m1_16911_22102# m1_16452_21590# m1_16452_21590# pfet$198
Xpfet$198_15 vdd m1_354_22513# m1_354_22513# m1_n46_22402# m1_488_21786# m1_488_21786#
+ pfet$198
Xnfet$228_1 m1_30256_19792# vss m1_32818_20470# vss nfet$228
Xnfet$235_2 m1_n6788_16080# m1_n6788_16080# m1_n7247_17714# m1_n7247_17714# m1_n6690_16398#
+ vss nfet$235
Xnfet$214_7 m1_n7383_17599# m1_n7383_17599# vss vss m1_n63_20470# vss nfet$214
Xnfet$216_17 m1_25107_21786# vss m1_25739_21786# vss nfet$216
Xnfet$232_16 m1_25722_20152# m1_25722_20152# m1_n3206_20274# m1_n3206_20274# m1_24556_20470#
+ vss nfet$232
Xpfet$225_0 vdd m1_n6380_21786# m1_n6380_21786# m1_n5019_19550# m1_n5227_20152# m1_n5227_20152#
+ pfet$225
Xnfet$240_0 m1_n9952_24224# m1_n9952_24224# m1_n10308_24542# m1_n10308_24542# m1_n9854_24542#
+ vss nfet$240
Xpfet$204_12 vdd vdd m1_32193_25858# m1_25107_21786# pfet$204
Xpfet$204_5 vdd vdd m1_326_24346# m1_n7513_20152# pfet$204
Xnfet$212_4 m1_2912_25858# vss m1_3049_25662# vss nfet$212
Xpfet$196_92 vdd vdd m1_28492_25858# m1_29607_24346# pfet$196
Xpfet$196_81 vdd vdd m1_18339_24542# m1_15943_25858# pfet$196
Xpfet$196_70 vdd vdd m1_14156_24542# m1_11760_25858# pfet$196
Xpfet$202_2 vdd vdd m1_1103_20152# m1_n7401_15478# pfet$202
Xpfet$201_13 vdd vdd m1_25747_17714# m1_26217_17714# pfet$201
Xnfet$239_9 m1_n3184_24224# vss m1_n3541_23922# vss nfet$239
Xnfet$224_17 m1_29256_21786# m1_29256_21786# vss vss m1_28094_21586# vss nfet$224
Xpfet$198_27 vdd m1_14422_22513# m1_14422_22513# m1_14022_22402# m1_14556_21786# m1_14556_21786#
+ pfet$198
Xpfet$198_16 vdd m1_24973_22513# m1_24973_22513# m1_23945_22102# m1_25739_21786# m1_25739_21786#
+ pfet$198
Xnfet$228_2 m1_31535_19792# m1_32818_20470# vss vss nfet$228
Xnfet$235_3 m1_n6172_16202# m1_n6172_16202# vss vss m1_n6690_16398# vss nfet$235
Xnfet$214_8 m1_27003_19550# m1_27003_19550# vss vss m1_27441_20470# vss nfet$214
Xnfet$232_17 m1_21880_15478# m1_21880_15478# m1_n3206_20274# m1_n3206_20274# m1_23924_20470#
+ vss nfet$232
Xnfet$233_0 m1_35837_22102# vss m1_n7513_20152# vss nfet$233
Xnfet$240_1 m1_n9336_24346# m1_n9336_24346# m1_n8625_26174# m1_n8625_26174# m1_n8389_25502#
+ vss nfet$240
Xpfet$225_1 vdd vdd vdd m1_n5019_22344# m1_n4485_21904# m1_n4485_21904# pfet$225
Xpfet$218_0 vdd m1_n10309_25662# m1_n10572_23922# m1_n10796_25662# pfet$218
Xpfet$204_13 vdd vdd m1_33790_24346# m1_n7513_20152# pfet$204
Xnfet$212_5 m1_2912_25858# m1_3536_25662# m1_3273_23922# vss nfet$212
Xpfet$204_6 vdd vdd m1_n290_24224# m1_n910_23922# pfet$204
Xpfet$196_93 vdd m1_28991_24224# m1_30095_25658# m1_28010_25858# pfet$196
Xpfet$196_82 vdd vdd m1_21241_24346# m1_n7513_20152# pfet$196
Xpfet$196_71 vdd vdd m1_11039_21786# m1_11760_25858# pfet$196
Xpfet$196_60 vdd vdd m1_20126_25858# m1_21241_24346# pfet$196
Xpfet$202_3 vdd vdd m1_5901_19550# m1_649_17714# pfet$202
Xpfet$200_0 vdd vdd m1_n1133_21590# m1_n1263_21786# pfet$200
Xpfet$198_28 vdd m1_14422_22513# m1_14422_22513# m1_13394_22102# m1_15188_21786# m1_15188_21786#
+ pfet$198
Xpfet$198_17 vdd m1_21456_22513# m1_21456_22513# m1_21056_22402# m1_21590_21786# m1_21590_21786#
+ pfet$198
Xnfet$235_4 m1_28113_15778# m1_28113_15778# m1_28003_18030# m1_28003_18030# m1_28239_17358#
+ vss nfet$235
Xnfet$228_3 m1_30256_22102# vss m1_32818_21586# vss nfet$228
Xnfet$214_9 m1_25747_17714# m1_25747_17714# vss vss m1_28073_20470# vss nfet$214
Xpfet$198_0 vdd vdd vdd m1_n674_22102# m1_n1133_21590# m1_n1133_21590# pfet$198
Xnfet$226_0 m1_34843_21786# m1_34843_21786# m1_34093_22102# m1_34093_22102# m1_34329_21430#
+ vss nfet$226
Xnfet$240_2 m1_n8848_25658# m1_n8848_25658# vss vss m1_n8389_25502# vss nfet$240
Xpfet$225_2 vdd m1_n5764_21786# m1_n5764_21786# m1_n5019_22344# m1_n5227_21418# m1_n5227_21418#
+ pfet$225
Xpfet$218_1 vdd m1_n9952_24224# m1_n8848_25658# m1_n10933_25858# pfet$218
Xnfet$212_6 m1_3049_25662# m1_3893_24224# m1_4997_25658# vss nfet$212
Xpfet$204_7 vdd vdd m1_32330_25662# m1_32193_25858# pfet$204
Xpfet$196_94 vdd m1_28492_25858# vdd m1_30095_25658# pfet$196
Xpfet$196_83 vdd m1_21729_25658# m1_22522_24542# m1_19781_25662# pfet$196
Xpfet$196_72 vdd m1_13363_25658# m1_14156_24542# m1_11415_25662# pfet$196
Xpfet$196_61 vdd m1_24452_24542# vdd m1_25424_24346# pfet$196
Xpfet$196_50 vdd vdd m1_20268_25662# m1_20126_25858# pfet$196
Xpfet$202_4 vdd vdd m1_12935_19550# m1_9015_17714# pfet$202
Xpfet$200_1 vdd vdd m1_11671_21786# m1_11039_21786# pfet$200
Xpfet$198_29 vdd vdd vdd m1_14022_22402# m1_12805_21786# m1_12805_21786# pfet$198
Xpfet$198_18 vdd vdd vdd m1_24573_22402# m1_23356_21786# m1_23356_21786# pfet$198
Xnfet$235_5 m1_26676_16080# m1_26676_16080# vss vss m1_28239_17358# vss nfet$235
Xnfet$211_20 m1_21241_24346# m1_21241_24346# m1_20126_25858# m1_20126_25858# m1_22188_25502#
+ vss nfet$211
Xpfet$198_1 vdd m1_7388_22513# m1_7388_22513# m1_6988_22402# m1_7522_21786# m1_7522_21786#
+ pfet$198
Xnfet$226_1 m1_28490_22513# m1_28490_22513# vss vss m1_34329_21430# vss nfet$226
Xnfet$219_0 m1_n3534_17714# vss m1_n6433_17343# vss nfet$219
Xnfet$240_3 m1_n9336_24346# m1_n9336_24346# vss vss m1_n9854_24542# vss nfet$240
Xpfet$218_2 vdd m1_n4362_24346# m1_n4847_25662# m1_n4464_25980# pfet$218
Xnfet$212_7 m1_3049_25662# m1_3273_23922# m1_3537_24542# vss nfet$212
Xpfet$204_8 vdd vdd m1_33174_24224# m1_32554_23922# pfet$204
Xpfet$196_95 vdd vdd m1_28991_24224# m1_28371_23922# pfet$196
Xpfet$196_84 vdd vdd m1_23827_25858# m1_18073_21786# pfet$196
Xpfet$196_73 vdd m1_16086_24542# vdd m1_17058_24346# pfet$196
Xpfet$196_62 vdd vdd m1_24452_24542# m1_24808_24224# pfet$196
Xpfet$196_51 vdd vdd m1_20625_24224# m1_20005_23922# pfet$196
Xpfet$196_40 vdd vdd m1_11760_25858# m1_12875_24346# pfet$196
Xpfet$223_0 vdd vdd m1_n7186_25858# m1_n10452_25858# pfet$223
Xpfet$202_5 vdd vdd m1_8137_20152# m1_965_15478# pfet$202
Xpfet$200_2 vdd vdd m1_12935_21590# m1_12805_21786# pfet$200
Xpfet$198_19 vdd m1_24973_22513# m1_24973_22513# m1_24573_22402# m1_25107_21786# m1_25107_21786#
+ pfet$198
Xnfet$235_6 m1_27292_16202# m1_27292_16202# vss vss m1_26774_16398# vss nfet$235
Xnfet$211_21 m1_28991_24224# m1_28991_24224# m1_28635_24542# m1_28635_24542# m1_29089_24542#
+ vss nfet$211
Xnfet$211_10 m1_17546_25658# m1_17546_25658# vss vss m1_18005_25502# vss nfet$211
Xpfet$198_2 vdd m1_7388_22513# m1_7388_22513# m1_6360_22102# m1_8154_21786# m1_8154_21786#
+ pfet$198
Xnfet$240_4 m1_n4978_24224# m1_n4978_24224# m1_n10452_25858# m1_n10452_25858# m1_n4880_24542#
+ vss nfet$240
Xnfet$226_2 m1_9645_21447# m1_9645_21447# vss vss m1_30492_21430# vss nfet$226
Xnfet$219_1 m1_n7513_20152# vss m1_n6788_16080# vss nfet$219
Xpfet$218_3 vdd m1_n3184_24224# m1_n3651_26174# m1_n4623_25487# pfet$218
Xnfet$212_8 m1_3394_25858# vss m1_3536_25662# vss nfet$212
Xpfet$204_9 vdd vdd m1_28624_21786# m1_32675_25947# pfet$204
Xnfet$231_0 m1_7198_15778# m1_7198_15778# m1_7088_18030# m1_7088_18030# m1_7324_17358#
+ vss nfet$231
Xpfet$196_41 vdd vdd m1_9288_21786# pd4 pfet$196
Xpfet$216_0 vdd vdd m1_n7513_20152# m1_35837_22102# pfet$216
Xpfet$196_30 vdd vdd m1_2912_25858# m1_488_21786# pfet$196
Xpfet$223_1 vdd m1_n7186_25858# vdd m1_n6111_25858# pfet$223
Xpfet$196_96 vdd m1_28635_24542# vdd m1_29607_24346# pfet$196
Xpfet$196_85 vdd m1_24188_23922# m1_24452_24542# m1_23827_25858# pfet$196
Xpfet$196_74 vdd vdd m1_14556_21786# m1_15943_25858# pfet$196
Xpfet$196_63 vdd vdd m1_19781_25662# m1_19644_25858# pfet$196
Xpfet$196_52 vdd m1_20268_25662# m1_20005_23922# m1_19781_25662# pfet$196
Xpfet$202_6 vdd vdd m1_9418_19550# m1_4832_17714# pfet$202
Xpfet$200_3 vdd vdd m1_9418_21590# m1_9288_21786# pfet$200
Xnfet$214_10 m1_9015_17714# m1_9015_17714# vss vss m1_14005_20470# vss nfet$214
Xnfet$235_7 m1_26676_16080# m1_26676_16080# m1_26217_17714# m1_26217_17714# m1_26774_16398#
+ vss nfet$235
Xnfet$211_22 m1_29607_24346# m1_29607_24346# vss vss m1_29089_24542# vss nfet$211
Xnfet$211_11 m1_16442_24224# m1_16442_24224# m1_16086_24542# m1_16086_24542# m1_16540_24542#
+ vss nfet$211
Xpfet$198_3 vdd m1_9645_21447# m1_9645_21447# m1_10505_22402# m1_11039_21786# m1_11039_21786#
+ pfet$198
Xpfet$199_30 vdd vdd vdd m1_24560_19550# m1_21880_15478# m1_21880_15478# pfet$199
Xnfet$226_3 m1_7388_22513# m1_7388_22513# m1_30256_22102# m1_30256_22102# m1_30492_21430#
+ vss nfet$226
Xnfet$219_2 m1_n4994_16080# vss m1_n5351_15778# vss nfet$219
Xnfet$240_5 m1_n4362_24346# m1_n4362_24346# vss vss m1_n4880_24542# vss nfet$240
Xpfet$218_4 vdd m1_n2567_23922# m1_n3184_24224# m1_n4464_25980# pfet$218
Xpfet$196_0 vdd vdd m1_3049_25662# m1_2912_25858# pfet$196
Xnfet$212_9 m1_3273_23922# vss m1_3893_24224# vss nfet$212
Xnfet$231_1 m1_5761_16080# m1_5761_16080# vss vss m1_7324_17358# vss nfet$231
Xnfet$224_0 m1_11039_21786# m1_11039_21786# vss vss m1_9877_21586# vss nfet$224
Xnfet$217_10 m1_26063_15478# vss m1_29239_20152# vss nfet$217
Xpfet$209_0 vdd vdd m1_n1263_21786# pd1 pfet$209
Xpfet$196_97 vdd vdd m1_21590_21786# m1_24309_25858# pfet$196
Xpfet$196_86 vdd m1_28634_25662# m1_28371_23922# m1_28147_25662# pfet$196
Xpfet$196_75 vdd vdd m1_19644_25858# m1_14556_21786# pfet$196
Xpfet$196_64 vdd vdd m1_22522_24542# m1_20126_25858# pfet$196
Xpfet$196_53 vdd m1_20625_24224# m1_21729_25658# m1_19644_25858# pfet$196
Xpfet$196_42 vdd m1_11760_25858# vdd m1_13363_25658# pfet$196
Xpfet$196_31 vdd m1_3273_23922# m1_3537_24542# m1_2912_25858# pfet$196
Xpfet$196_20 vdd vdd m1_4509_24346# m1_n7513_20152# pfet$196
Xpfet$202_7 vdd vdd m1_11654_20152# m1_5148_15478# pfet$202
Xnfet$214_11 m1_13198_17714# m1_13198_17714# vss vss m1_17522_20470# vss nfet$214
Xpfet$200_4 vdd vdd m1_8154_21786# m1_7522_21786# pfet$200
Xpfet$198_4 vdd vdd vdd m1_9877_22102# m1_9418_21590# m1_9418_21590# pfet$198
Xnfet$211_23 m1_25424_24346# m1_25424_24346# m1_24309_25858# m1_24309_25858# m1_26371_25502#
+ vss nfet$211
Xnfet$211_12 m1_17058_24346# m1_17058_24346# m1_15943_25858# m1_15943_25858# m1_18005_25502#
+ vss nfet$211
Xpfet$199_31 vdd m1_n2543_20130# m1_n2543_20130# m1_20407_19850# m1_19969_19550# m1_19969_19550#
+ pfet$199
Xpfet$199_20 vdd m1_n3822_21786# m1_n3822_21786# m1_14009_19550# m1_9015_17714# m1_9015_17714#
+ pfet$199
Xnfet$219_3 m1_n6433_17343# vss m1_n6274_17836# vss nfet$219
Xnfet$240_6 m1_n4978_24224# m1_n4978_24224# vss vss m1_n3415_25502# vss nfet$240
Xpfet$196_1 vdd m1_3536_25662# m1_3273_23922# m1_3049_25662# pfet$196
Xpfet$218_5 vdd m1_n10572_23922# m1_n10308_24542# m1_n10933_25858# pfet$218
Xpfet$209_1 vdd vdd m1_2254_21786# pd2 pfet$209
Xnfet$217_0 m1_n3534_17714# vss m1_2384_19550# vss nfet$217
Xnfet$231_2 m1_9944_16080# m1_9944_16080# vss vss m1_11507_17358# vss nfet$231
Xnfet$224_1 m1_11671_21786# m1_11671_21786# vss vss m1_10509_21586# vss nfet$224
Xpfet$196_98 vdd m1_30095_25658# m1_30888_24542# m1_28147_25662# pfet$196
Xpfet$196_87 vdd vdd m1_28147_25662# m1_28010_25858# pfet$196
Xpfet$196_76 vdd m1_20005_23922# m1_20269_24542# m1_19644_25858# pfet$196
Xpfet$196_65 vdd vdd m1_18073_21786# m1_20126_25858# pfet$196
Xpfet$196_54 vdd vdd m1_24808_24224# m1_24188_23922# pfet$196
Xpfet$196_43 vdd vdd m1_12805_21786# pd5 pfet$196
Xnfet$217_11 m1_9331_15478# vss m1_15171_20152# vss nfet$217
Xpfet$196_32 vdd vdd m1_7720_24542# m1_8076_24224# pfet$196
Xpfet$196_21 vdd m1_7456_23922# m1_7720_24542# m1_7095_25858# pfet$196
Xpfet$196_10 vdd m1_8076_24224# m1_9180_25658# m1_7095_25858# pfet$196
Xpfet$202_8 vdd vdd m1_n1133_19550# m1_n7383_17599# pfet$202
Xpfet$221_0 vdd vdd m1_n4485_20152# m1_n3822_20130# pfet$221
Xnfet$214_12 m1_16452_19550# m1_16452_19550# vss vss m1_16890_20470# vss nfet$214
Xpfet$200_5 vdd vdd m1_1120_21786# m1_488_21786# pfet$200
Xnfet$247_0 m1_n6839_20152# vss m1_n8145_21908# vss nfet$247
Xnfet$211_24 m1_30095_25658# m1_30095_25658# vss vss m1_30554_25502# vss nfet$211
Xnfet$211_13 m1_13363_25658# m1_13363_25658# vss vss m1_13822_25502# vss nfet$211
Xpfet$199_32 vdd m1_n2543_20130# m1_n2543_20130# m1_21043_19550# m1_17381_17714# m1_17381_17714#
+ pfet$199
Xpfet$199_21 vdd vdd vdd m1_13373_19850# m1_15171_20152# m1_15171_20152# pfet$199
Xpfet$199_10 vdd vdd vdd m1_9856_19850# m1_11654_20152# m1_11654_20152# pfet$199
Xpfet$198_5 vdd m1_9645_21447# m1_9645_21447# m1_9877_22102# m1_11671_21786# m1_11671_21786#
+ pfet$198
Xnfet$219_4 m1_n7247_17714# vss m1_n4377_15778# vss nfet$219
Xnfet$240_7 m1_n3541_23922# m1_n3541_23922# m1_n3651_26174# m1_n3651_26174# m1_n3415_25502#
+ vss nfet$240
Xpfet$196_2 vdd vdd m1_3394_25858# m1_4509_24346# pfet$196
Xpfet$218_6 vdd m1_n8848_25658# m1_n8055_24542# m1_n10796_25662# pfet$218
Xnfet$217_1 m1_n3218_15478# vss m1_4620_20152# vss nfet$217
Xnfet$231_3 m1_11381_15778# m1_11381_15778# m1_11271_18030# m1_11271_18030# m1_11507_17358#
+ vss nfet$231
Xnfet$224_2 m1_8154_21786# m1_8154_21786# vss vss m1_6992_21586# vss nfet$224
Xpfet$196_99 vdd vdd m1_26705_24542# m1_24309_25858# pfet$196
Xpfet$209_2 vdd vdd m1_26873_21786# pd9 pfet$209
Xpfet$196_88 vdd vdd m1_28634_25662# m1_28492_25858# pfet$196
Xpfet$196_77 vdd vdd m1_20269_24542# m1_20625_24224# pfet$196
Xpfet$196_66 vdd vdd m1_15461_25858# m1_11039_21786# pfet$196
Xpfet$196_55 vdd m1_24451_25662# m1_24188_23922# m1_23964_25662# pfet$196
Xpfet$196_44 vdd m1_15943_25858# vdd m1_17546_25658# pfet$196
Xnfet$217_12 m1_13514_15478# vss m1_18688_20152# vss nfet$217
Xpfet$196_33 vdd vdd m1_7522_21786# m1_7577_25858# pfet$196
Xpfet$196_22 vdd vdd m1_3537_24542# m1_3893_24224# pfet$196
Xpfet$196_11 vdd vdd m1_7719_25662# m1_7577_25858# pfet$196
Xpfet$202_9 vdd vdd m1_27003_19550# m1_25747_17714# pfet$202
Xpfet$214_0 vdd vdd m1_n7247_17714# m1_n6788_16080# pfet$214
Xpfet$221_1 vdd m1_n4485_21904# vdd m1_9624_19404# pfet$221
Xnfet$214_13 m1_19969_19550# m1_19969_19550# vss vss m1_20407_20470# vss nfet$214
Xpfet$200_6 vdd vdd m1_5901_21590# m1_5771_21786# pfet$200
Xnfet$239_10 vss vss m1_n4978_24224# vss nfet$239
Xnfet$211_25 m1_29607_24346# m1_29607_24346# m1_28492_25858# m1_28492_25858# m1_30554_25502#
+ vss nfet$211
Xnfet$211_14 m1_12875_24346# m1_12875_24346# m1_11760_25858# m1_11760_25858# m1_13822_25502#
+ vss nfet$211
Xpfet$198_6 vdd vdd vdd m1_10505_22402# m1_9288_21786# m1_9288_21786# pfet$198
Xpfet$199_33 vdd m1_n3206_20274# m1_n3206_20274# m1_24560_19550# m1_21564_17714# m1_21564_17714#
+ pfet$199
Xpfet$199_22 vdd vdd vdd m1_14009_19550# m1_9331_15478# m1_9331_15478# pfet$199
Xpfet$199_11 vdd vdd vdd m1_10492_19550# m1_5148_15478# m1_5148_15478# pfet$199
Xnfet$219_5 m1_n7247_17714# vss m1_n6657_17518# vss nfet$219
Xpfet$196_3 vdd m1_3394_25858# vdd m1_4997_25658# pfet$196
Xpfet$218_7 vdd m1_n3541_23922# m1_n4362_24346# m1_n4623_25487# pfet$218
Xnfet$217_2 m1_n7401_15478# vss m1_1103_20152# vss nfet$217
Xnfet$231_4 m1_10560_16202# m1_10560_16202# vss vss m1_10042_16398# vss nfet$231
Xnfet$224_3 m1_7522_21786# m1_7522_21786# vss vss m1_6360_21586# vss nfet$224
Xpfet$196_89 vdd vdd m1_19839_21786# pd7 pfet$196
Xpfet$196_78 vdd m1_20269_24542# vdd m1_21241_24346# pfet$196
Xpfet$196_67 vdd m1_15822_23922# m1_16086_24542# m1_15461_25858# pfet$196
Xpfet$196_56 vdd m1_24808_24224# m1_25912_25658# m1_23827_25858# pfet$196
Xpfet$196_45 vdd vdd m1_16442_24224# m1_15822_23922# pfet$196
Xnfet$217_13 m1_13198_17714# vss m1_16452_19550# vss nfet$217
Xpfet$196_34 vdd m1_9180_25658# m1_9973_24542# m1_7232_25662# pfet$196
Xpfet$196_23 vdd m1_3537_24542# vdd m1_4509_24346# pfet$196
Xpfet$196_12 vdd m1_7577_25858# vdd m1_9180_25658# pfet$196
Xpfet$207_0 vdd m1_31535_19792# vdd m1_17939_22513# pfet$207
Xnfet$222_0 pd1 vss m1_n1263_21786# vss nfet$222
Xpfet$214_1 vdd m1_n7247_17714# vdd m1_n6172_16202# pfet$214
Xpfet$221_2 vdd m1_n5227_21418# vdd m1_2590_19404# pfet$221
Xpfet$200_7 vdd vdd m1_4637_21786# m1_4005_21786# pfet$200
Xnfet$214_14 m1_17381_17714# m1_17381_17714# vss vss m1_21039_20470# vss nfet$214
Xnfet$239_11 m1_n10452_25858# vss m1_n4847_25662# vss nfet$239
Xpfet$197_110 vdd vdd m1_10458_17836# m1_10299_17343# pfet$197
Xnfet$211_26 m1_25912_25658# m1_25912_25658# vss vss m1_26371_25502# vss nfet$211
Xnfet$211_15 m1_25424_24346# m1_25424_24346# vss vss m1_24906_24542# vss nfet$211
Xpfet$198_7 vdd m1_354_22513# m1_354_22513# m1_n674_22102# m1_1120_21786# m1_1120_21786#
+ pfet$198
Xpfet$199_34 vdd m1_n3206_20274# m1_n3206_20274# m1_23924_19850# m1_23486_19550# m1_23486_19550#
+ pfet$199
Xpfet$199_23 vdd vdd vdd m1_16890_19850# m1_18688_20152# m1_18688_20152# pfet$199
Xpfet$199_12 vdd m1_6107_19404# m1_6107_19404# m1_6975_19550# m1_649_17714# m1_649_17714#
+ pfet$199
Xnfet$219_6 m1_n7247_17714# vss m1_n7383_17599# vss nfet$219
Xpfet$196_4 vdd vdd m1_3893_24224# m1_3273_23922# pfet$196
Xnfet$212_80 m1_28147_25662# m1_28991_24224# m1_30095_25658# vss nfet$212
Xnfet$217_3 m1_649_17714# vss m1_5901_19550# vss nfet$217
Xnfet$231_5 m1_9944_16080# m1_9944_16080# m1_9485_17714# m1_9485_17714# m1_10042_16398#
+ vss nfet$231
Xnfet$224_4 m1_1120_21786# m1_1120_21786# vss vss m1_n42_21586# vss nfet$224
Xpfet$196_57 vdd vdd m1_24451_25662# m1_24309_25858# pfet$196
Xpfet$196_46 vdd m1_16442_24224# m1_17546_25658# m1_15461_25858# pfet$196
Xnfet$217_14 m1_21564_17714# vss m1_23486_19550# vss nfet$217
Xpfet$196_35 vdd m1_7720_24542# vdd m1_8692_24346# pfet$196
Xpfet$196_24 vdd vdd m1_5790_24542# m1_3394_25858# pfet$196
Xpfet$196_13 vdd vdd m1_12259_24224# m1_11639_23922# pfet$196
Xpfet$196_79 vdd m1_17546_25658# m1_18339_24542# m1_15598_25662# pfet$196
Xpfet$196_68 vdd vdd m1_16086_24542# m1_16442_24224# pfet$196
Xnfet$222_1 pd2 vss m1_2254_21786# vss nfet$222
Xnfet$215_0 m1_9485_17714# vss m1_9015_17714# vss nfet$215
Xpfet$207_1 vdd vdd m1_30256_19792# m1_21456_22513# pfet$207
Xpfet$214_2 vdd vdd m1_n5461_18030# m1_n5351_15778# pfet$214
Xpfet$221_3 vdd vdd m1_n5227_21418# m1_6107_19404# pfet$221
Xpfet$200_8 vdd vdd m1_2384_21590# m1_2254_21786# pfet$200
Xnfet$214_15 m1_21564_17714# m1_21564_17714# vss vss m1_24556_20470# vss nfet$214
Xnfet$239_12 m1_n10452_25858# vss m1_n5571_25662# vss nfet$239
Xpfet$202_10 vdd vdd m1_29239_20152# m1_26063_15478# pfet$202
Xpfet$197_100 vdd vdd m1_23820_18030# m1_23930_15778# pfet$197
Xnfet$215_80 m1_18824_17836# m1_19747_15778# m1_18926_16202# vss nfet$215
Xnfet$211_27 m1_12875_24346# m1_12875_24346# vss vss m1_12357_24542# vss nfet$211
Xnfet$211_16 m1_24808_24224# m1_24808_24224# m1_24452_24542# m1_24452_24542# m1_24906_24542#
+ vss nfet$211
Xpfet$198_8 vdd vdd vdd m1_6360_22102# m1_5901_21590# m1_5901_21590# pfet$198
Xpfet$199_35 vdd m1_n3822_21786# m1_n3822_21786# m1_13373_19850# m1_12935_19550# m1_12935_19550#
+ pfet$199
Xpfet$199_24 vdd m1_n1927_20274# m1_n1927_20274# m1_16890_19850# m1_16452_19550# m1_16452_19550#
+ pfet$199
Xpfet$199_13 vdd m1_n927_19404# m1_n927_19404# m1_n695_19850# m1_n1133_19550# m1_n1133_19550#
+ pfet$199
Xnfet$219_7 m1_26217_17714# vss m1_26807_17518# vss nfet$219
Xnfet$245_0 m1_n927_19404# m1_n927_19404# vss vss m1_n6282_20470# vss nfet$245
Xpfet$196_5 vdd m1_3893_24224# m1_4997_25658# m1_2912_25858# pfet$196
Xnfet$212_81 m1_n7513_20152# vss m1_25424_24346# vss nfet$212
Xnfet$212_70 m1_21590_21786# vss m1_28010_25858# vss nfet$212
Xnfet$217_4 m1_4832_17714# vss m1_9418_19550# vss nfet$217
Xnfet$231_6 m1_1578_16080# m1_1578_16080# vss vss m1_3141_17358# vss nfet$231
Xnfet$224_5 m1_4005_21786# m1_4005_21786# vss vss m1_2843_21586# vss nfet$224
Xnfet$217_15 m1_17697_15478# vss m1_22205_20152# vss nfet$217
Xpfet$196_69 vdd vdd m1_12875_24346# m1_n7513_20152# pfet$196
Xpfet$196_58 vdd vdd m1_23964_25662# m1_23827_25858# pfet$196
Xpfet$196_47 vdd vdd m1_15943_25858# m1_17058_24346# pfet$196
Xpfet$196_36 vdd vdd m1_8692_24346# m1_n7513_20152# pfet$196
Xpfet$196_25 vdd vdd m1_4005_21786# m1_3394_25858# pfet$196
Xpfet$196_14 vdd vdd m1_11902_25662# m1_11760_25858# pfet$196
Xnfet$222_2 pd9 vss m1_26873_21786# vss nfet$222
Xnfet$215_1 m1_9015_17714# vss m1_6116_17343# vss nfet$215
Xpfet$207_2 vdd m1_30256_19792# vdd m1_24973_22513# pfet$207
Xpfet$214_3 vdd m1_n5461_18030# vdd m1_n6788_16080# pfet$214
Xpfet$221_4 vdd vdd m1_n4485_21904# m1_n3822_21786# pfet$221
Xpfet$197_90 vdd m1_19747_15778# m1_18926_16202# m1_18665_17343# pfet$197
Xpfet$212_0 vdd vdd fout m1_34093_22102# pfet$212
Xpfet$200_9 vdd vdd m1_22222_21786# m1_21590_21786# pfet$200
Xnfet$214_16 m1_23486_19550# m1_23486_19550# vss vss m1_23924_20470# vss nfet$214
Xnfet$239_13 fin vss m1_n4623_25487# vss nfet$239
Xpfet$197_101 vdd vdd m1_19637_18030# m1_19747_15778# pfet$197
Xpfet$202_11 vdd vdd m1_18688_20152# m1_13514_15478# pfet$202
Xnfet$215_81 m1_13198_17714# vss m1_10299_17343# vss nfet$215
Xnfet$215_70 m1_n7513_20152# vss m1_18310_16080# vss nfet$215
Xpfet$198_9 vdd m1_3871_22513# m1_3871_22513# m1_3471_22402# m1_4005_21786# m1_4005_21786#
+ pfet$198
Xnfet$211_17 m1_20625_24224# m1_20625_24224# m1_20269_24542# m1_20269_24542# m1_20723_24542#
+ vss nfet$211
Xpfet$199_25 vdd vdd vdd m1_17526_19550# m1_13514_15478# m1_13514_15478# pfet$199
Xpfet$199_14 vdd m1_n927_19404# m1_n927_19404# m1_n59_19550# m1_n7383_17599# m1_n7383_17599#
+ pfet$199
Xnfet$219_8 m1_n7513_20152# vss m1_26676_16080# vss nfet$219
Xpfet$196_6 vdd vdd m1_3536_25662# m1_3394_25858# pfet$196
Xnfet$238_0 m1_n3822_20130# m1_n3822_20130# m1_n4485_20152# m1_n4485_20152# m1_n3724_20470#
+ vss nfet$238
Xnfet$245_1 m1_n2543_20130# m1_n2543_20130# m1_n5227_20152# m1_n5227_20152# m1_n2445_20470#
+ vss nfet$245
Xnfet$212_82 m1_11415_25662# m1_12259_24224# m1_13363_25658# vss nfet$212
Xnfet$212_71 m1_28147_25662# m1_28371_23922# m1_28635_24542# vss nfet$212
Xnfet$212_60 pd6 vss m1_16322_21786# vss nfet$212
Xnfet$217_5 m1_965_15478# vss m1_8137_20152# vss nfet$217
Xnfet$231_7 m1_5761_16080# m1_5761_16080# m1_5302_17714# m1_5302_17714# m1_5859_16398#
+ vss nfet$231
Xnfet$224_6 m1_4637_21786# m1_4637_21786# vss vss m1_3475_21586# vss nfet$224
Xpfet$196_59 vdd vdd m1_16322_21786# pd6 pfet$196
Xpfet$196_48 vdd m1_16085_25662# m1_15822_23922# m1_15598_25662# pfet$196
Xnfet$217_16 m1_17381_17714# vss m1_19969_19550# vss nfet$217
Xpfet$196_37 vdd vdd m1_9973_24542# m1_7577_25858# pfet$196
Xpfet$196_26 vdd m1_4997_25658# m1_5790_24542# m1_3049_25662# pfet$196
Xpfet$196_15 vdd m1_11902_25662# m1_11639_23922# m1_11415_25662# pfet$196
Xnfet$215_2 m1_6275_17836# m1_7555_16080# m1_7088_18030# vss nfet$215
Xpfet$207_3 vdd vdd m1_34843_21786# m1_34093_19792# pfet$207
Xpfet$214_4 vdd vdd m1_26217_17714# m1_26676_16080# pfet$214
Xpfet$221_5 vdd m1_n6839_21786# vdd m1_n5764_21786# pfet$221
Xpfet$197_91 vdd m1_24287_16080# m1_23820_18030# m1_22848_17343# pfet$197
Xpfet$197_80 vdd vdd m1_15564_15778# m1_15921_16080# pfet$197
Xnfet$214_17 m1_12935_19550# m1_12935_19550# vss vss m1_13373_20470# vss nfet$214
Xnfet$220_0 m1_n10452_25858# vss m1_n1271_25858# vss nfet$220
Xpfet$205_0 vdd vdd m1_n646_24542# m1_n290_24224# pfet$205
Xpfet$202_12 vdd vdd m1_15171_20152# m1_9331_15478# pfet$202
Xpfet$197_102 vdd vdd m1_13198_17714# m1_13668_17714# pfet$197
Xnfet$215_82 m1_10299_17343# vss m1_10458_17836# vss nfet$215
Xnfet$215_71 m1_14641_17836# m1_15921_16080# m1_15454_18030# vss nfet$215
Xnfet$215_60 m1_18665_17343# vss m1_18824_17836# vss nfet$215
Xnfet$211_18 m1_21241_24346# m1_21241_24346# vss vss m1_20723_24542# vss nfet$211
Xpfet$199_26 vdd m1_n1927_20274# m1_n1927_20274# m1_17526_19550# m1_13198_17714# m1_13198_17714#
+ pfet$199
Xpfet$199_15 vdd vdd vdd m1_n59_19550# m1_n7401_15478# m1_n7401_15478# pfet$199
Xnfet$219_9 m1_n10452_25858# vss m1_27031_17343# vss nfet$219
.ends

.subckt pfet$265 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$263 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$283 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt nfet$281 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$264 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$262 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$284 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$282 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt asc_drive_buffer vss in vdd out
Xpfet$265_0 vdd vdd m1_3466_n454# in pfet$265
Xpfet$263_0 m1_4274_n1060# vdd vdd m1_4274_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ vdd m1_4002_n1060# m1_4002_n1060# pfet$263
Xnfet$283_0 m1_3466_n454# vss m1_4002_n1060# vss nfet$283
Xnfet$281_0 m1_4274_n1060# vss m1_4002_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ m1_4274_n1060# vss m1_4002_n1060# vss nfet$281
Xpfet$264_0 vdd vdd m1_4002_n1060# m1_3466_n454# pfet$264
Xpfet$262_0 out out m1_4274_n1060# vdd m1_4274_n1060# out vdd vdd m1_4274_n1060# out
+ m1_4274_n1060# m1_4274_n1060# out m1_4274_n1060# vdd m1_4274_n1060# vdd m1_4274_n1060#
+ pfet$262
Xnfet$284_0 in vss m1_3466_n454# vss nfet$284
Xnfet$282_0 out out vss m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# m1_4274_n1060#
+ m1_4274_n1060# out m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# vss vss
+ nfet$282
.ends

.subckt pfet$244 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$242 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$268 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$273 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$240 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$266 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$259 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$271 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$264 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$249 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$254 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$262 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$247 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$252 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$245 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$260 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$250 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$243 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$269 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$241 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$267 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$272 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$265 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$270 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$263 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$248 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$253 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$246 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$261 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$251 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt asc_lock_detector_20250826 ref vdd div lock vss
Xpfet$244_4 vdd vdd m1_15618_394# m1_12790_n340# pfet$244
Xpfet$242_1 m1_12790_n340# m1_12790_n340# m1_11642_n340# vdd m1_11642_n340# m1_12790_n340#
+ vdd vdd m1_11642_n340# m1_12790_n340# m1_11642_n340# m1_11642_n340# m1_12790_n340#
+ m1_11642_n340# vdd m1_11642_n340# vdd m1_11642_n340# pfet$242
Xnfet$268_1 m1_15618_394# vss m1_15755_n208# vss nfet$268
Xpfet$244_5 vdd vdd m1_17215_2028# vss pfet$244
Xpfet$242_2 m1_4402_n340# m1_4402_n340# m1_3254_n340# vdd m1_3254_n340# m1_4402_n340#
+ vdd vdd m1_3254_n340# m1_4402_n340# m1_3254_n340# m1_3254_n340# m1_4402_n340# m1_3254_n340#
+ vdd m1_3254_n340# vdd m1_3254_n340# pfet$242
Xnfet$268_2 m1_n2336_5099# vss m1_16242_n208# vss nfet$268
Xnfet$273_0 m1_19675_2344# vss lock vss nfet$273
Xpfet$244_6 vdd vdd m1_19469_1832# m1_17926_34# pfet$244
Xpfet$240_0 vdd vdd m1_6640_1478# m1_4402_n340# pfet$240
Xpfet$242_3 m1_208_n340# m1_208_n340# m1_n940_n340# vdd m1_n940_n340# m1_208_n340#
+ vdd vdd m1_n940_n340# m1_208_n340# m1_n940_n340# m1_n940_n340# m1_208_n340# m1_n940_n340#
+ vdd m1_n940_n340# vdd m1_n940_n340# pfet$242
Xnfet$268_3 m1_17926_34# vss m1_18496_1828# vss nfet$268
Xnfet$266_0 m1_15755_n208# m1_16599_2028# m1_17703_788# vss nfet$266
Xpfet$244_7 vdd vdd m1_17215_5644# vss pfet$244
Xpfet$242_4 m1_208_7868# m1_208_7868# m1_n940_4493# vdd m1_n940_4493# m1_208_7868#
+ vdd vdd m1_n940_4493# m1_208_7868# m1_n940_4493# m1_n940_4493# m1_208_7868# m1_n940_4493#
+ vdd m1_n940_4493# vdd m1_n940_4493# pfet$242
Xpfet$240_1 vdd vdd m1_10834_1478# m1_8596_n340# pfet$240
Xnfet$266_1 m1_15618_394# m1_16242_n208# m1_15979_2344# vss nfet$266
Xnfet$259_0 m1_8596_n340# m1_8596_n340# vss m1_7448_n340# m1_7448_n340# m1_8596_n340#
+ vss m1_7448_n340# m1_7448_n340# m1_7448_n340# m1_8596_n340# m1_7448_n340# m1_7448_n340#
+ m1_8596_n340# vss m1_7448_n340# vss vss nfet$259
Xnfet$268_4 m1_12790_n340# vss m1_15618_394# vss nfet$268
Xpfet$244_8 vdd vdd m1_19469_4920# m1_17926_7472# pfet$244
Xpfet$242_5 m1_12790_7868# m1_12790_7868# m1_11642_4493# vdd m1_11642_4493# m1_12790_7868#
+ vdd vdd m1_11642_4493# m1_12790_7868# m1_11642_4493# m1_11642_4493# m1_12790_7868#
+ m1_11642_4493# vdd m1_11642_4493# vdd m1_11642_4493# pfet$242
Xpfet$240_2 vdd vdd m1_n1748_1478# ref pfet$240
Xnfet$268_5 vss vss m1_17215_2028# vss nfet$268
Xnfet$259_1 m1_4402_n340# m1_4402_n340# vss m1_3254_n340# m1_3254_n340# m1_4402_n340#
+ vss m1_3254_n340# m1_3254_n340# m1_3254_n340# m1_4402_n340# m1_3254_n340# m1_3254_n340#
+ m1_4402_n340# vss m1_3254_n340# vss vss nfet$259
Xnfet$266_2 m1_15618_394# m1_17703_788# m1_18496_1828# vss nfet$266
Xpfet$242_6 m1_4402_7868# m1_4402_7868# m1_3254_4493# vdd m1_3254_4493# m1_4402_7868#
+ vdd vdd m1_3254_4493# m1_4402_7868# m1_3254_4493# m1_3254_4493# m1_4402_7868# m1_3254_4493#
+ vdd m1_3254_4493# vdd m1_3254_4493# pfet$242
Xpfet$244_9 vdd vdd m1_18496_5840# m1_17926_7472# pfet$244
Xnfet$271_0 m1_n4030_5270# vss m1_n2336_5099# vss nfet$271
Xpfet$240_3 vdd vdd m1_n1748_5099# m1_n2336_5099# pfet$240
Xnfet$259_2 m1_12790_n340# m1_12790_n340# vss m1_11642_n340# m1_11642_n340# m1_12790_n340#
+ vss m1_11642_n340# m1_11642_n340# m1_11642_n340# m1_12790_n340# m1_11642_n340# m1_11642_n340#
+ m1_12790_n340# vss m1_11642_n340# vss vss nfet$259
Xnfet$266_3 m1_15755_n208# m1_15979_2344# m1_16243_1828# vss nfet$266
Xnfet$268_6 m1_17926_34# vss m1_19469_1832# vss nfet$268
Xnfet$264_0 m1_n7214_4493# vss m1_n7486_4493# m1_n7486_4493# m1_n7486_4493# m1_n7214_4493#
+ m1_n7214_4493# vss m1_n7486_4493# vss nfet$264
Xpfet$249_0 vdd vdd m1_n11680_4493# m1_n12216_5099# pfet$249
Xpfet$242_7 m1_8596_7868# m1_8596_7868# m1_7448_4493# vdd m1_7448_4493# m1_8596_7868#
+ vdd vdd m1_7448_4493# m1_8596_7868# m1_7448_4493# m1_7448_4493# m1_8596_7868# m1_7448_4493#
+ vdd m1_7448_4493# vdd m1_7448_4493# pfet$242
Xpfet$240_4 vdd vdd m1_6640_5099# m1_4402_7868# pfet$240
Xnfet$268_7 vss vss m1_17215_5644# vss nfet$268
Xnfet$266_4 m1_15618_7156# m1_17703_6956# m1_18496_5840# vss nfet$266
Xnfet$259_3 m1_208_n340# m1_208_n340# vss m1_n940_n340# m1_n940_n340# m1_208_n340#
+ vss m1_n940_n340# m1_n940_n340# m1_n940_n340# m1_208_n340# m1_n940_n340# m1_n940_n340#
+ m1_208_n340# vss m1_n940_n340# vss vss nfet$259
Xnfet$264_1 m1_n15602_4493# vss m1_n15874_4493# m1_n15874_4493# m1_n15874_4493# m1_n15602_4493#
+ m1_n15602_4493# vss m1_n15874_4493# vss nfet$264
Xpfet$249_1 vdd vdd m1_n7486_4493# m1_n8022_5099# pfet$249
Xpfet$240_5 vdd vdd m1_10834_5099# m1_8596_7868# pfet$240
Xnfet$268_8 m1_17926_7472# vss m1_19469_4920# vss nfet$268
Xnfet$259_4 m1_12790_7868# m1_12790_7868# vss m1_11642_4493# m1_11642_4493# m1_12790_7868#
+ vss m1_11642_4493# m1_11642_4493# m1_11642_4493# m1_12790_7868# m1_11642_4493# m1_11642_4493#
+ m1_12790_7868# vss m1_11642_4493# vss vss nfet$259
Xnfet$264_2 m1_n11408_4493# vss m1_n11680_4493# m1_n11680_4493# m1_n11680_4493# m1_n11408_4493#
+ m1_n11408_4493# vss m1_n11680_4493# vss nfet$264
Xnfet$266_5 m1_15755_6960# m1_15979_5220# m1_16243_5840# vss nfet$266
Xpfet$249_2 vdd vdd m1_n15874_4493# m1_n16410_5099# pfet$249
Xpfet$240_6 vdd vdd m1_2446_5099# m1_208_7868# pfet$240
Xpfet$254_0 vdd vdd lock m1_19675_2344# pfet$254
Xnfet$268_9 m1_17926_7472# vss m1_18496_5840# vss nfet$268
Xnfet$259_5 m1_8596_7868# m1_8596_7868# vss m1_7448_4493# m1_7448_4493# m1_8596_7868#
+ vss m1_7448_4493# m1_7448_4493# m1_7448_4493# m1_8596_7868# m1_7448_4493# m1_7448_4493#
+ m1_8596_7868# vss m1_7448_4493# vss vss nfet$259
Xnfet$266_6 m1_15618_7156# m1_16242_6960# m1_15979_5220# vss nfet$266
Xnfet$262_0 m1_n6066_7868# m1_n6066_7868# vss m1_n7214_4493# m1_n7214_4493# m1_n6066_7868#
+ vss m1_n7214_4493# m1_n7214_4493# m1_n7214_4493# m1_n6066_7868# m1_n7214_4493# m1_n7214_4493#
+ m1_n6066_7868# vss m1_n7214_4493# vss vss nfet$262
Xpfet$240_7 vdd vdd m1_2446_1478# m1_208_n340# pfet$240
Xpfet$247_0 m1_n10260_7868# m1_n10260_7868# m1_n11408_4493# vdd m1_n11408_4493# m1_n10260_7868#
+ vdd vdd m1_n11408_4493# m1_n10260_7868# m1_n11408_4493# m1_n11408_4493# m1_n10260_7868#
+ m1_n11408_4493# vdd m1_n11408_4493# vdd m1_n11408_4493# pfet$247
Xnfet$259_6 m1_208_7868# m1_208_7868# vss m1_n940_4493# m1_n940_4493# m1_208_7868#
+ vss m1_n940_4493# m1_n940_4493# m1_n940_4493# m1_208_7868# m1_n940_4493# m1_n940_4493#
+ m1_208_7868# vss m1_n940_4493# vss vss nfet$259
Xnfet$266_7 m1_15755_6960# m1_16599_5522# m1_17703_6956# vss nfet$266
Xnfet$262_1 m1_n14454_7868# m1_n14454_7868# vss m1_n15602_4493# m1_n15602_4493# m1_n14454_7868#
+ vss m1_n15602_4493# m1_n15602_4493# m1_n15602_4493# m1_n14454_7868# m1_n15602_4493#
+ m1_n15602_4493# m1_n14454_7868# vss m1_n15602_4493# vss vss nfet$262
Xpfet$247_1 m1_n6066_7868# m1_n6066_7868# m1_n7214_4493# vdd m1_n7214_4493# m1_n6066_7868#
+ vdd vdd m1_n7214_4493# m1_n6066_7868# m1_n7214_4493# m1_n7214_4493# m1_n6066_7868#
+ m1_n7214_4493# vdd m1_n7214_4493# vdd m1_n7214_4493# pfet$247
Xnfet$259_7 m1_4402_7868# m1_4402_7868# vss m1_3254_4493# m1_3254_4493# m1_4402_7868#
+ vss m1_3254_4493# m1_3254_4493# m1_3254_4493# m1_4402_7868# m1_3254_4493# m1_3254_4493#
+ m1_4402_7868# vss m1_3254_4493# vss vss nfet$259
Xnfet$262_2 m1_n10260_7868# m1_n10260_7868# vss m1_n11408_4493# m1_n11408_4493# m1_n10260_7868#
+ vss m1_n11408_4493# m1_n11408_4493# m1_n11408_4493# m1_n10260_7868# m1_n11408_4493#
+ m1_n11408_4493# m1_n10260_7868# vss m1_n11408_4493# vss vss nfet$262
Xpfet$252_0 vdd vdd m1_n2336_5099# m1_n4030_5270# pfet$252
Xpfet$247_2 m1_n14454_7868# m1_n14454_7868# m1_n15602_4493# vdd m1_n15602_4493# m1_n14454_7868#
+ vdd vdd m1_n15602_4493# m1_n14454_7868# m1_n15602_4493# m1_n15602_4493# m1_n14454_7868#
+ m1_n15602_4493# vdd m1_n15602_4493# vdd m1_n15602_4493# pfet$247
Xpfet$245_0 vdd m1_16599_2028# m1_17703_788# m1_15618_394# pfet$245
Xnfet$260_0 m1_10834_1478# vss m1_11370_n340# vss nfet$260
Xpfet$245_1 vdd m1_16242_n208# m1_15979_2344# m1_15755_n208# pfet$245
Xnfet$260_1 m1_2446_1478# vss m1_2982_n340# vss nfet$260
Xpfet$244_10 vdd vdd m1_15618_7156# m1_12790_7868# pfet$244
Xnfet$260_2 m1_6640_1478# vss m1_7176_n340# vss nfet$260
Xpfet$245_2 vdd m1_15979_2344# m1_16243_1828# m1_15618_394# pfet$245
Xpfet$250_0 vdd vdd m1_n8022_5099# m1_n10260_7868# pfet$250
Xpfet$244_11 vdd vdd m1_16599_5522# m1_15979_5220# pfet$244
Xnfet$260_3 m1_n1748_1478# vss m1_n1212_n340# vss nfet$260
Xpfet$245_3 vdd m1_17703_788# m1_18496_1828# m1_15755_n208# pfet$245
Xpfet$243_0 m1_7448_n340# vdd vdd m1_7448_n340# m1_7176_n340# m1_7176_n340# m1_7448_n340#
+ vdd m1_7176_n340# m1_7176_n340# pfet$243
Xpfet$250_1 vdd vdd m1_n16410_5099# div pfet$250
Xpfet$244_12 vdd vdd m1_16242_6960# ref pfet$244
Xnfet$269_0 m1_n14454_7868# vss m1_n12216_5099# vss nfet$269
Xnfet$260_4 m1_10834_5099# vss m1_11370_4493# vss nfet$260
Xpfet$245_4 vdd m1_17703_6956# m1_18496_5840# m1_15755_6960# pfet$245
Xpfet$243_1 m1_11642_n340# vdd vdd m1_11642_n340# m1_11370_n340# m1_11370_n340# m1_11642_n340#
+ vdd m1_11370_n340# m1_11370_n340# pfet$243
Xpfet$250_2 vdd vdd m1_n12216_5099# m1_n14454_7868# pfet$250
Xpfet$244_13 vdd vdd m1_15755_6960# m1_15618_7156# pfet$244
Xnfet$269_1 div vss m1_n16410_5099# vss nfet$269
Xnfet$260_5 m1_6640_5099# vss m1_7176_4493# vss nfet$260
Xpfet$245_5 vdd m1_15979_5220# m1_16243_5840# m1_15618_7156# pfet$245
Xpfet$243_2 m1_3254_n340# vdd vdd m1_3254_n340# m1_2982_n340# m1_2982_n340# m1_3254_n340#
+ vdd m1_2982_n340# m1_2982_n340# pfet$243
Xnfet$269_2 m1_n10260_7868# vss m1_n8022_5099# vss nfet$269
Xnfet$260_6 m1_n1748_5099# vss m1_n1212_4493# vss nfet$260
Xpfet$245_6 vdd m1_16599_5522# m1_17703_6956# m1_15618_7156# pfet$245
Xpfet$243_3 m1_n940_n340# vdd vdd m1_n940_n340# m1_n1212_n340# m1_n1212_n340# m1_n940_n340#
+ vdd m1_n1212_n340# m1_n1212_n340# pfet$243
Xpfet$241_0 vdd vdd m1_7176_n340# m1_6640_1478# pfet$241
Xnfet$267_0 m1_17215_2028# m1_17215_2028# m1_17926_34# m1_17926_34# m1_18162_712#
+ vss nfet$267
Xnfet$260_7 m1_2446_5099# vss m1_2982_4493# vss nfet$260
Xpfet$245_7 vdd m1_16242_6960# m1_15979_5220# m1_15755_6960# pfet$245
Xpfet$243_4 m1_n940_4493# vdd vdd m1_n940_4493# m1_n1212_4493# m1_n1212_4493# m1_n940_4493#
+ vdd m1_n1212_4493# m1_n1212_4493# pfet$243
Xpfet$241_1 vdd vdd m1_11370_n340# m1_10834_1478# pfet$241
Xnfet$267_1 m1_17703_788# m1_17703_788# vss vss m1_18162_712# vss nfet$267
Xpfet$243_5 m1_11642_4493# vdd vdd m1_11642_4493# m1_11370_4493# m1_11370_4493# m1_11642_4493#
+ vdd m1_11370_4493# m1_11370_4493# pfet$243
Xpfet$241_2 vdd vdd m1_2982_n340# m1_2446_1478# pfet$241
Xnfet$267_2 m1_16599_2028# m1_16599_2028# m1_16243_1828# m1_16243_1828# m1_16697_1672#
+ vss nfet$267
Xnfet$272_0 m1_19469_4920# m1_19469_4920# m1_19675_2344# m1_19675_2344# m1_19911_1672#
+ vss nfet$272
Xpfet$243_6 m1_3254_4493# vdd vdd m1_3254_4493# m1_2982_4493# m1_2982_4493# m1_3254_4493#
+ vdd m1_2982_4493# m1_2982_4493# pfet$243
Xpfet$241_3 vdd vdd m1_n1212_n340# m1_n1748_1478# pfet$241
Xnfet$268_10 m1_12790_7868# vss m1_15618_7156# vss nfet$268
Xnfet$265_0 m1_8596_n340# vss m1_10834_1478# vss nfet$265
Xnfet$267_3 m1_17215_2028# m1_17215_2028# vss vss m1_16697_1672# vss nfet$267
Xnfet$272_1 m1_19469_1832# m1_19469_1832# vss vss m1_19911_1672# vss nfet$272
Xpfet$243_7 m1_7448_4493# vdd vdd m1_7448_4493# m1_7176_4493# m1_7176_4493# m1_7448_4493#
+ vdd m1_7176_4493# m1_7176_4493# pfet$243
Xpfet$241_4 vdd vdd m1_n1212_4493# m1_n1748_5099# pfet$241
Xnfet$268_11 m1_15979_5220# vss m1_16599_5522# vss nfet$268
Xnfet$267_4 m1_17215_5644# m1_17215_5644# vss vss m1_16697_5840# vss nfet$267
Xnfet$265_1 m1_4402_n340# vss m1_6640_1478# vss nfet$265
Xpfet$241_5 vdd vdd m1_2982_4493# m1_2446_5099# pfet$241
Xnfet$268_12 m1_15618_7156# vss m1_15755_6960# vss nfet$268
Xnfet$267_5 m1_16599_5522# m1_16599_5522# m1_16243_5840# m1_16243_5840# m1_16697_5840#
+ vss nfet$267
Xnfet$265_2 ref vss m1_n1748_1478# vss nfet$265
Xnfet$270_0 div m1_n4030_5270# vss vss nfet$270
Xpfet$241_6 vdd vdd m1_7176_4493# m1_6640_5099# pfet$241
Xnfet$267_6 m1_17215_5644# m1_17215_5644# m1_17926_7472# m1_17926_7472# m1_18162_6800#
+ vss nfet$267
Xnfet$268_13 ref vss m1_16242_6960# vss nfet$268
Xnfet$265_3 m1_n2336_5099# vss m1_n1748_5099# vss nfet$265
Xnfet$263_0 m1_n8022_5099# vss m1_n7486_4493# vss nfet$263
Xpfet$241_7 vdd vdd m1_11370_4493# m1_10834_5099# pfet$241
Xnfet$270_1 m1_n6066_7868# vss m1_n4030_5270# vss nfet$270
Xpfet$248_0 m1_n11408_4493# vdd vdd m1_n11408_4493# m1_n11680_4493# m1_n11680_4493#
+ m1_n11408_4493# vdd m1_n11680_4493# m1_n11680_4493# pfet$248
Xnfet$267_7 m1_17703_6956# m1_17703_6956# vss vss m1_18162_6800# vss nfet$267
Xnfet$263_1 m1_n16410_5099# vss m1_n15874_4493# vss nfet$263
Xnfet$265_4 m1_8596_7868# vss m1_10834_5099# vss nfet$265
Xpfet$248_1 m1_n7214_4493# vdd vdd m1_n7214_4493# m1_n7486_4493# m1_n7486_4493# m1_n7214_4493#
+ vdd m1_n7486_4493# m1_n7486_4493# pfet$248
Xnfet$265_5 m1_4402_7868# vss m1_6640_5099# vss nfet$265
Xnfet$263_2 m1_n12216_5099# vss m1_n11680_4493# vss nfet$263
Xpfet$248_2 m1_n15602_4493# vdd vdd m1_n15602_4493# m1_n15874_4493# m1_n15874_4493#
+ m1_n15602_4493# vdd m1_n15874_4493# m1_n15874_4493# pfet$248
Xpfet$253_0 vdd m1_19675_2344# vdd m1_19469_1832# pfet$253
Xnfet$265_6 m1_208_n340# vss m1_2446_1478# vss nfet$265
Xpfet$246_0 vdd m1_17926_34# vdd m1_17703_788# pfet$246
Xnfet$261_0 m1_3254_n340# vss m1_2982_n340# m1_2982_n340# m1_2982_n340# m1_3254_n340#
+ m1_3254_n340# vss m1_2982_n340# vss nfet$261
Xpfet$253_1 vdd vdd m1_19675_2344# m1_19469_4920# pfet$253
Xnfet$265_7 m1_208_7868# vss m1_2446_5099# vss nfet$265
Xpfet$246_1 vdd vdd m1_17926_34# m1_17215_2028# pfet$246
Xnfet$261_1 m1_7448_n340# vss m1_7176_n340# m1_7176_n340# m1_7176_n340# m1_7448_n340#
+ m1_7448_n340# vss m1_7176_n340# vss nfet$261
Xpfet$246_2 vdd m1_16243_1828# vdd m1_17215_2028# pfet$246
Xnfet$261_2 m1_11642_n340# vss m1_11370_n340# m1_11370_n340# m1_11370_n340# m1_11642_n340#
+ m1_11642_n340# vss m1_11370_n340# vss nfet$261
Xpfet$251_0 vdd vdd vdd m1_n3798_6028# div div pfet$251
Xpfet$246_3 vdd vdd m1_16243_1828# m1_16599_2028# pfet$246
Xnfet$261_3 m1_n940_n340# vss m1_n1212_n340# m1_n1212_n340# m1_n1212_n340# m1_n940_n340#
+ m1_n940_n340# vss m1_n1212_n340# vss nfet$261
Xpfet$244_0 vdd vdd m1_16599_2028# m1_15979_2344# pfet$244
Xpfet$251_1 vdd m1_n4030_5270# m1_n4030_5270# m1_n3798_6028# m1_n6066_7868# m1_n6066_7868#
+ pfet$251
Xnfet$261_4 m1_11642_4493# vss m1_11370_4493# m1_11370_4493# m1_11370_4493# m1_11642_4493#
+ m1_11642_4493# vss m1_11370_4493# vss nfet$261
Xpfet$246_4 vdd m1_16243_5840# vdd m1_17215_5644# pfet$246
Xpfet$244_1 vdd vdd m1_16242_n208# m1_n2336_5099# pfet$244
Xnfet$261_5 m1_7448_4493# vss m1_7176_4493# m1_7176_4493# m1_7176_4493# m1_7448_4493#
+ m1_7448_4493# vss m1_7176_4493# vss nfet$261
Xpfet$246_5 vdd vdd m1_16243_5840# m1_16599_5522# pfet$246
Xpfet$244_2 vdd vdd m1_15755_n208# m1_15618_394# pfet$244
Xnfet$261_6 m1_n940_4493# vss m1_n1212_4493# m1_n1212_4493# m1_n1212_4493# m1_n940_4493#
+ m1_n940_4493# vss m1_n1212_4493# vss nfet$261
Xpfet$246_6 vdd m1_17926_7472# vdd m1_17703_6956# pfet$246
Xpfet$244_3 vdd vdd m1_18496_1828# m1_17926_34# pfet$244
Xpfet$242_0 m1_8596_n340# m1_8596_n340# m1_7448_n340# vdd m1_7448_n340# m1_8596_n340#
+ vdd vdd m1_7448_n340# m1_8596_n340# m1_7448_n340# m1_7448_n340# m1_8596_n340# m1_7448_n340#
+ vdd m1_7448_n340# vdd m1_7448_n340# pfet$242
Xnfet$268_0 m1_15979_2344# vss m1_16599_2028# vss nfet$268
Xnfet$261_7 m1_3254_4493# vss m1_2982_4493# m1_2982_4493# m1_2982_4493# m1_3254_4493#
+ m1_3254_4493# vss m1_2982_4493# vss nfet$261
Xpfet$246_7 vdd vdd m1_17926_7472# m1_17215_5644# pfet$246
.ends

.subckt pfet$256 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$274 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$255 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$275 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt xp_3_1_MUX S0 S1 VDD VSS OUT_1 C_1 B_1 A_1
Xpfet$256_0 VDD VDD m1_n432_n1290# S1 pfet$256
Xpfet$256_1 VDD VDD m1_n432_458# S0 pfet$256
Xnfet$274_0 m1_n432_n1290# C_1 OUT_1 VSS nfet$274
Xnfet$274_1 m1_n432_458# B_1 m1_239_n318# VSS nfet$274
Xnfet$274_3 S0 A_1 m1_239_n318# VSS nfet$274
Xnfet$274_2 S1 m1_239_n318# OUT_1 VSS nfet$274
Xpfet$255_0 VDD A_1 m1_239_n318# m1_n432_458# pfet$255
Xpfet$255_1 VDD C_1 OUT_1 S1 pfet$255
Xpfet$255_2 VDD B_1 m1_239_n318# S0 pfet$255
Xpfet$255_3 VDD m1_239_n318# OUT_1 m1_n432_n1290# pfet$255
Xnfet$275_0 S1 VSS m1_n432_n1290# VSS nfet$275
Xnfet$275_1 S0 VSS m1_n432_458# VSS nfet$275
.ends

.subckt nfet$250 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt nfet$249 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$233 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$252 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt inv1u05u VDD in VSS out
Xpfet$233_0 VDD VDD out in pfet$233
Xnfet$252_0 in VSS out VSS nfet$252
.ends

.subckt pfet$231 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=4.55p ps=15.3u w=7u l=0.5u
.ends

.subckt nfet$248 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt nfet$251 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$232 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pass1u05u VDD VSS ind ins clkp clkn
Xnfet$251_0 clkn ind ins VSS nfet$251
Xpfet$232_0 VDD ind ins clkp pfet$232
.ends

.subckt nfet$253 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$229 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_954_0# w_n180_n88# a_854_n136#
+ a_n92_0# a_446_n136# a_650_n136# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt pfet$234 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.5u
.ends

.subckt pfet$230 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_954_0# w_n180_n88#
+ a_38_n60# a_n92_0# a_1058_n60# a_854_n60# a_342_0# a_138_0# a_650_n60#
X0 a_954_0# a_854_n60# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n60# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt xp_programmable_basic_pump up vdd s1 s2 s3 s4 down out iref vss
Xnfet$250_0 m1_n7879_n12170# pass1u05u_0/ins m1_n7879_n12170# out pass1u05u_0/ins
+ vss nfet$250
Xnfet$249_9 down down vss vss m1_n8807_n11192# vss nfet$249
Xinv1u05u_3 vdd s1 vss inv1u05u_3/out inv1u05u
Xnfet$250_1 m1_n7879_n12170# pass1u05u_0/ins m1_n7879_n12170# out pass1u05u_0/ins
+ vss nfet$250
Xnfet$250_2 vss down vss m1_n7879_n12170# down vss nfet$250
Xnfet$250_3 vss down vss m1_n7879_n12170# down vss nfet$250
Xnfet$250_4 vss down vss m1_n7879_n12170# down vss nfet$250
Xnfet$250_5 vss down vss m1_n7879_n12170# down vss nfet$250
Xnfet$250_6 m1_n7879_n12170# pass1u05u_0/ins m1_n7879_n12170# out pass1u05u_0/ins
+ vss nfet$250
Xpfet$231_0 vdd vdd vdd vdd pfet$231
Xnfet$250_7 m1_n7879_n12170# pass1u05u_0/ins m1_n7879_n12170# out pass1u05u_0/ins
+ vss nfet$250
Xnfet$250_10 m1_n8607_n8040# pass1u05u_1/ins m1_n8607_n8040# out pass1u05u_1/ins vss
+ nfet$250
Xpfet$231_1 vdd vdd vdd vdd pfet$231
Xnfet$250_8 vss vdd vss m1_n8144_n9165# vdd vss nfet$250
Xnfet$248_10 pass1u05u_2/ins pass1u05u_2/ins m1_n7679_n8960# m1_n7679_n8960# out vss
+ nfet$248
Xnfet$250_11 m1_n8144_n9165# iref m1_n8144_n9165# iref iref vss nfet$250
Xpfet$231_2 vdd vdd vdd vdd pfet$231
Xnfet$250_9 m1_n7216_n8262# iref m1_n7216_n8262# pass1u05u_7/ind iref vss nfet$250
Xnfet$248_11 vss vss vss vss vss vss nfet$248
Xnfet$250_12 vss down vss m1_n8607_n8040# down vss nfet$250
Xpfet$231_3 vdd vdd vdd vdd pfet$231
Xnfet$248_12 down down vss vss m1_n7679_n8960# vss nfet$248
Xnfet$250_13 vss vdd vss m1_n7216_n8262# vdd vss nfet$250
Xpfet$231_4 vdd vdd vdd vdd pfet$231
Xpass1u05u_0 vdd vss iref pass1u05u_0/ins inv1u05u_1/out s3 pass1u05u
Xnfet$248_13 vss vss vss vss vss vss nfet$248
Xnfet$248_0 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$248
Xnfet$250_14 m1_n8607_n8040# pass1u05u_1/ins m1_n8607_n8040# out pass1u05u_1/ins vss
+ nfet$250
Xpfet$231_5 vdd vdd vdd vdd pfet$231
Xpass1u05u_1 vdd vss iref pass1u05u_1/ins inv1u05u_2/out s2 pass1u05u
Xnfet$248_14 vss vss vss vss vss vss nfet$248
Xnfet$248_1 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$248
Xnfet$250_15 vss down vss m1_n8607_n8040# down vss nfet$250
Xpfet$231_6 vdd vdd vdd vdd pfet$231
Xpass1u05u_2 vdd vss iref pass1u05u_2/ins inv1u05u_3/out s1 pass1u05u
Xnfet$248_15 vss vss vss vss vss vss nfet$248
Xnfet$253_0 inv1u05u_2/out pass1u05u_1/ins vss vss nfet$253
Xnfet$248_2 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$248
Xpfet$231_7 vdd vdd vdd vdd pfet$231
Xpass1u05u_3 vdd vss pass1u05u_7/ind pass1u05u_3/ins inv1u05u_3/out s1 pass1u05u
Xnfet$248_3 vss vss vss vss vss vss nfet$248
Xnfet$253_1 inv1u05u_3/out pass1u05u_2/ins vss vss nfet$253
Xpfet$231_8 vdd vdd vdd vdd pfet$231
Xpass1u05u_4 vdd vss pass1u05u_7/ind pass1u05u_4/ins inv1u05u_2/out s2 pass1u05u
Xnfet$253_2 inv1u05u_0/out pass1u05u_6/ins vss vss nfet$253
Xnfet$248_4 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$248
Xpfet$231_9 vdd vdd vdd vdd pfet$231
Xpass1u05u_5 vdd vss pass1u05u_7/ind pass1u05u_5/ins inv1u05u_1/out s3 pass1u05u
Xnfet$248_5 vss vss vss vss vss vss nfet$248
Xnfet$253_3 inv1u05u_1/out pass1u05u_0/ins vss vss nfet$253
Xpass1u05u_6 vdd vss iref pass1u05u_6/ins inv1u05u_0/out s4 pass1u05u
Xnfet$248_6 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$248
Xpfet$229_0 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$229
Xpass1u05u_7 vdd vss pass1u05u_7/ind pass1u05u_7/ins inv1u05u_0/out s4 pass1u05u
Xnfet$248_7 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$248
Xpfet$229_1 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$229
Xnfet$248_8 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$248
Xpfet$229_2 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$229
Xpfet$234_0 vdd s3 pass1u05u_5/ins vdd pfet$234
Xnfet$248_9 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$248
Xnfet$249_10 vss vss vss vss vss vss nfet$249
Xpfet$229_3 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$229
Xpfet$234_1 vdd s2 pass1u05u_4/ins vdd pfet$234
Xnfet$249_11 vss vss vss vss vss vss nfet$249
Xpfet$234_2 vdd s1 pass1u05u_3/ins vdd pfet$234
Xpfet$229_4 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$229
Xnfet$249_12 vss vss vss vss vss vss nfet$249
Xpfet$229_5 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$229
Xpfet$234_3 vdd s4 pass1u05u_7/ins vdd pfet$234
Xpfet$231_20 vdd vdd vdd vdd pfet$231
Xnfet$249_13 vss vss vss vss vss vss nfet$249
Xpfet$229_6 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$229
Xpfet$229_20 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$229
Xpfet$231_21 vdd vdd vdd vdd pfet$231
Xpfet$231_10 vdd vdd vdd vdd pfet$231
Xpfet$229_7 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$229
Xpfet$229_21 m1_n6703_2564# m1_n6703_2564# pass1u05u_4/ins out out vdd pass1u05u_4/ins
+ m1_n6703_2564# pass1u05u_4/ins pass1u05u_4/ins m1_n6703_2564# out pass1u05u_4/ins
+ pass1u05u_4/ins pfet$229
Xpfet$231_22 vdd vdd vdd vdd pfet$231
Xpfet$229_10 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$229
Xpfet$231_11 vdd vdd vdd vdd pfet$231
Xpfet$229_8 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$229
Xpfet$229_22 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$229
Xpfet$229_11 vdd vdd up m1_n5450_4559# m1_n5450_4559# vdd up vdd up up vdd m1_n5450_4559#
+ up up pfet$229
Xpfet$231_23 vdd vdd vdd vdd pfet$231
Xpfet$230_0 vdd vdd m1_n4127_3649# vss vss m1_n4127_3649# vdd vss vdd vss vss vdd
+ m1_n4127_3649# vss pfet$230
Xpfet$231_12 vdd vdd vdd vdd pfet$231
Xpfet$229_9 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$229
Xpfet$229_23 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$229
Xpfet$229_12 vdd vdd up m1_n6703_2564# m1_n6703_2564# vdd up vdd up up vdd m1_n6703_2564#
+ up up pfet$229
Xpfet$230_1 m1_n5580_883# m1_n5580_883# out pass1u05u_5/ins pass1u05u_5/ins out vdd
+ pass1u05u_5/ins m1_n5580_883# pass1u05u_5/ins pass1u05u_5/ins m1_n5580_883# out
+ pass1u05u_5/ins pfet$230
Xpfet$231_13 vdd vdd vdd vdd pfet$231
Xnfet$249_0 down down vss vss m1_n8807_n11192# vss nfet$249
Xpfet$229_24 m1_n5450_4559# m1_n5450_4559# pass1u05u_3/ins out out vdd pass1u05u_3/ins
+ m1_n5450_4559# pass1u05u_3/ins pass1u05u_3/ins m1_n5450_4559# out pass1u05u_3/ins
+ pass1u05u_3/ins pfet$229
Xpfet$231_14 vdd vdd vdd vdd pfet$231
Xpfet$229_13 vdd vdd up m1_n6703_2564# m1_n6703_2564# vdd up vdd up up vdd m1_n6703_2564#
+ up up pfet$229
Xpfet$230_2 m1_n5580_883# m1_n5580_883# out pass1u05u_5/ins pass1u05u_5/ins out vdd
+ pass1u05u_5/ins m1_n5580_883# pass1u05u_5/ins pass1u05u_5/ins m1_n5580_883# out
+ pass1u05u_5/ins pfet$230
Xnfet$249_1 down down vss vss m1_n8807_n11192# vss nfet$249
Xpfet$229_25 m1_n6703_2564# m1_n6703_2564# pass1u05u_4/ins out out vdd pass1u05u_4/ins
+ m1_n6703_2564# pass1u05u_4/ins pass1u05u_4/ins m1_n6703_2564# out pass1u05u_4/ins
+ pass1u05u_4/ins pfet$229
Xpfet$230_3 m1_n5580_883# m1_n5580_883# out pass1u05u_5/ins pass1u05u_5/ins out vdd
+ pass1u05u_5/ins m1_n5580_883# pass1u05u_5/ins pass1u05u_5/ins m1_n5580_883# out
+ pass1u05u_5/ins pfet$230
Xpfet$229_14 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$229
Xpfet$231_15 vdd vdd vdd vdd pfet$231
Xnfet$249_2 down down vss vss m1_n8807_n11192# vss nfet$249
Xpfet$231_16 vdd vdd vdd vdd pfet$231
Xpfet$230_4 m1_n5580_883# m1_n5580_883# out pass1u05u_5/ins pass1u05u_5/ins out vdd
+ pass1u05u_5/ins m1_n5580_883# pass1u05u_5/ins pass1u05u_5/ins m1_n5580_883# out
+ pass1u05u_5/ins pfet$230
Xpfet$229_15 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$229
Xnfet$249_3 down down vss vss m1_n8807_n11192# vss nfet$249
Xpfet$230_5 m1_n4127_3649# m1_n4127_3649# pass1u05u_7/ind pass1u05u_7/ind pass1u05u_7/ind
+ pass1u05u_7/ind vdd pass1u05u_7/ind m1_n4127_3649# pass1u05u_7/ind pass1u05u_7/ind
+ m1_n4127_3649# pass1u05u_7/ind pass1u05u_7/ind pfet$230
Xpfet$229_16 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$229
Xpfet$231_17 vdd vdd vdd vdd pfet$231
Xnfet$249_4 vss vss vss vss vss vss nfet$249
Xpfet$231_18 vdd vdd vdd vdd pfet$231
Xpfet$229_17 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$229
Xnfet$249_5 vss vss vss vss vss vss nfet$249
Xpfet$229_18 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$229
Xpfet$231_19 vdd vdd vdd vdd pfet$231
Xnfet$249_6 down down vss vss m1_n8807_n11192# vss nfet$249
Xinv1u05u_0 vdd s4 vss inv1u05u_0/out inv1u05u
Xpfet$229_19 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$229
Xnfet$249_7 down down vss vss m1_n8807_n11192# vss nfet$249
Xinv1u05u_1 vdd s3 vss inv1u05u_1/out inv1u05u
Xnfet$249_8 down down vss vss m1_n8807_n11192# vss nfet$249
Xinv1u05u_2 vdd s2 vss inv1u05u_2/out inv1u05u
.ends

.subckt pfet$235 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$257 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$255 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$238 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$236 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$258 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$256 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$254 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$239 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$237 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt asc_hysteresis_buffer$5 vss in vdd out
Xpfet$235_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd
+ m1_884_42# m1_884_42# pfet$235
Xnfet$257_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$257
Xnfet$255_0 m1_348_648# vss m1_884_42# vss nfet$255
Xpfet$238_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$238
Xpfet$236_0 vdd vdd m1_884_42# m1_348_648# pfet$236
Xnfet$258_0 m1_1156_42# vss m1_884_42# vss nfet$258
Xnfet$256_0 in vss m1_348_648# vss nfet$256
Xnfet$254_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$254
Xpfet$239_0 vdd vdd m1_884_42# m1_1156_42# pfet$239
Xpfet$237_0 vdd vdd m1_348_648# in pfet$237
.ends

.subckt xp_3_1_MUX$4 S0 S1 VDD VSS OUT_1 C_1 B_1 A_1
Xpfet$256_0 VDD VDD m1_n432_n1290# S1 pfet$256
Xpfet$256_1 VDD VDD m1_n432_458# S0 pfet$256
Xnfet$274_0 m1_n432_n1290# C_1 OUT_1 VSS nfet$274
Xnfet$274_1 m1_n432_458# B_1 m1_239_n318# VSS nfet$274
Xnfet$274_3 S0 A_1 m1_239_n318# VSS nfet$274
Xnfet$274_2 S1 m1_239_n318# OUT_1 VSS nfet$274
Xpfet$255_0 VDD A_1 m1_239_n318# m1_n432_458# pfet$255
Xpfet$255_1 VDD C_1 OUT_1 S1 pfet$255
Xpfet$255_2 VDD B_1 m1_239_n318# S0 pfet$255
Xpfet$255_3 VDD m1_239_n318# OUT_1 m1_n432_n1290# pfet$255
Xnfet$275_0 S1 VSS m1_n432_n1290# VSS nfet$275
Xnfet$275_1 S0 VSS m1_n432_458# VSS nfet$275
.ends

.subckt asc_dual_psd_def_20250809$4 vdd vss pd1 pd2 pd3 pd4 pd5 pd6 pd7 pd8 pd9 fout
+ sd1 sd2 sd3 sd4 sd5 sd6 sd7 sd8 sd9 fin define
Xpfet$196_7 vdd vdd m1_7232_25662# m1_7095_25858# pfet$196
Xnfet$238_1 m1_n1927_20274# m1_n1927_20274# vss vss m1_n2445_20470# vss nfet$238
Xnfet$212_72 m1_23827_25858# m1_25912_25658# m1_26705_24542# vss nfet$212
Xnfet$212_61 m1_23964_25662# m1_24808_24224# m1_25912_25658# vss nfet$212
Xnfet$212_50 m1_n7513_20152# vss m1_21241_24346# vss nfet$212
Xnfet$224_7 m1_488_21786# m1_488_21786# vss vss m1_n674_21586# vss nfet$224
Xnfet$217_6 m1_9015_17714# vss m1_12935_19550# vss nfet$217
Xnfet$231_8 m1_3015_15778# m1_3015_15778# m1_2905_18030# m1_2905_18030# m1_3141_17358#
+ vss nfet$231
Xnfet$217_17 m1_21880_15478# vss m1_25722_20152# vss nfet$217
Xpfet$196_49 vdd m1_20126_25858# vdd m1_21729_25658# pfet$196
Xpfet$196_38 vdd vdd m1_16085_25662# m1_15943_25858# pfet$196
Xpfet$196_27 vdd vdd m1_11278_25858# m1_7522_21786# pfet$196
Xpfet$196_16 vdd vdd m1_5771_21786# pd3 pfet$196
Xpfet$207_4 vdd m1_34093_19792# vdd m1_32818_20470# pfet$207
Xpfet$214_5 vdd m1_26217_17714# vdd m1_27292_16202# pfet$214
Xnfet$215_3 m1_n7513_20152# vss m1_9944_16080# vss nfet$215
Xpfet$221_6 vdd vdd m1_n6973_21481# m1_n6839_21786# pfet$221
Xpfet$197_92 vdd m1_15454_18030# vdd m1_14127_16080# pfet$197
Xpfet$197_81 vdd vdd m1_13668_17714# m1_14127_16080# pfet$197
Xpfet$197_70 vdd vdd m1_18824_17836# m1_18665_17343# pfet$197
Xnfet$213_0 m1_n1133_21590# m1_n1133_21590# m1_354_22513# m1_354_22513# m1_n674_21586#
+ vss nfet$213
Xnfet$220_1 m1_n789_25858# vss m1_n647_25662# vss nfet$220
Xpfet$205_1 vdd m1_n789_25858# vdd m1_814_25658# pfet$205
Xpfet$202_13 vdd vdd m1_16452_19550# m1_13198_17714# pfet$202
Xpfet$197_103 vdd m1_14743_16202# m1_14258_17518# m1_14641_17836# pfet$197
Xnfet$215_72 m1_17851_17714# vss m1_18441_17518# vss nfet$215
Xnfet$215_61 m1_20104_16080# vss m1_19747_15778# vss nfet$215
Xnfet$215_50 m1_25747_17714# vss m1_22848_17343# vss nfet$215
Xnfet$211_19 m1_21729_25658# m1_21729_25658# vss vss m1_22188_25502# vss nfet$211
Xpfet$199_27 vdd vdd vdd m1_20407_19850# m1_22205_20152# m1_22205_20152# pfet$199
Xpfet$199_16 vdd vdd vdd m1_28077_19550# m1_26063_15478# m1_26063_15478# pfet$199
Xpfet$196_8 vdd vdd m1_8076_24224# m1_7456_23922# pfet$196
Xnfet$238_2 m1_n3206_20274# m1_n3206_20274# vss vss m1_n3724_20470# vss nfet$238
Xnfet$212_73 m1_24309_25858# vss m1_21590_21786# vss nfet$212
Xnfet$212_62 m1_24188_23922# vss m1_24808_24224# vss nfet$212
Xnfet$212_51 m1_19644_25858# m1_21729_25658# m1_22522_24542# vss nfet$212
Xnfet$212_40 m1_15598_25662# m1_16442_24224# m1_17546_25658# vss nfet$212
Xnfet$224_8 m1_25739_21786# m1_25739_21786# vss vss m1_24577_21586# vss nfet$224
Xnfet$217_7 m1_5148_15478# vss m1_11654_20152# vss nfet$217
Xnfet$231_9 m1_2194_16202# m1_2194_16202# vss vss m1_1676_16398# vss nfet$231
Xpfet$196_39 vdd vdd m1_15598_25662# m1_15461_25858# pfet$196
Xpfet$196_28 vdd m1_11639_23922# m1_11903_24542# m1_11278_25858# pfet$196
Xpfet$196_17 vdd vdd m1_7577_25858# m1_8692_24346# pfet$196
Xnfet$243_0 m1_n8283_20611# vss m1_n8283_19850# vss nfet$243
Xpfet$228_0 vdd vdd m1_n8145_21908# m1_n6839_20152# pfet$228
Xpfet$214_6 vdd vdd m1_28003_18030# m1_28113_15778# pfet$214
Xpfet$207_5 vdd vdd m1_34093_19792# m1_32818_21586# pfet$207
Xnfet$215_4 m1_10299_17343# m1_10560_16202# m1_10075_17518# vss nfet$215
Xpfet$221_7 vdd vdd m1_n6839_21786# m1_n6380_21786# pfet$221
Xpfet$197_93 vdd m1_23820_18030# vdd m1_22493_16080# pfet$197
Xpfet$197_82 vdd m1_13668_17714# vdd m1_14743_16202# pfet$197
Xpfet$197_71 vdd vdd m1_19747_15778# m1_20104_16080# pfet$197
Xpfet$197_60 vdd vdd m1_n194_15778# m1_n3064_17714# pfet$197
Xnfet$213_1 m1_n1263_21786# m1_n1263_21786# m1_354_22513# m1_354_22513# m1_n42_21586#
+ vss nfet$213
Xnfet$220_2 m1_n1271_25858# vss m1_n1134_25662# vss nfet$220
Xpfet$205_2 vdd vdd m1_n789_25858# m1_326_24346# pfet$205
Xpfet$202_14 vdd vdd m1_23486_19550# m1_21564_17714# pfet$202
Xpfet$197_104 vdd vdd m1_14127_16080# m1_n7513_20152# pfet$197
Xpfet$210_0 vdd m1_34093_22102# vdd m1_28490_22513# pfet$210
Xnfet$215_73 m1_13668_17714# vss m1_16538_15778# vss nfet$215
Xnfet$215_62 m1_18665_17343# m1_20721_15778# m1_20104_16080# vss nfet$215
Xnfet$215_51 m1_n7513_20152# vss m1_22493_16080# vss nfet$215
Xnfet$215_40 m1_n2250_17343# m1_n194_15778# m1_n811_16080# vss nfet$215
Xpfet$199_28 vdd vdd vdd m1_21043_19550# m1_17697_15478# m1_17697_15478# pfet$199
Xpfet$199_17 vdd m1_n3822_20130# m1_n3822_20130# m1_28077_19550# m1_25747_17714# m1_25747_17714#
+ pfet$199
Xnfet$238_3 m1_n6973_21481# m1_n6973_21481# m1_n6839_20152# m1_n6839_20152# m1_n6282_20470#
+ vss nfet$238
Xpfet$196_9 vdd m1_7719_25662# m1_7456_23922# m1_7232_25662# pfet$196
Xnfet$212_74 pd8 vss m1_23356_21786# vss nfet$212
Xnfet$212_63 m1_14556_21786# vss m1_19644_25858# vss nfet$212
Xnfet$212_52 m1_20126_25858# vss m1_22522_24542# vss nfet$212
Xnfet$212_41 pd5 vss m1_12805_21786# vss nfet$212
Xnfet$212_30 m1_n7513_20152# vss m1_17058_24346# vss nfet$212
Xnfet$224_9 m1_25107_21786# m1_25107_21786# vss vss m1_23945_21586# vss nfet$224
Xnfet$217_8 m1_n7383_17599# vss m1_n1133_19550# vss nfet$217
Xpfet$196_29 vdd vdd m1_11903_24542# m1_12259_24224# pfet$196
Xpfet$196_18 vdd vdd m1_11415_25662# m1_11278_25858# pfet$196
Xnfet$243_1 m1_n7513_20152# m1_n8283_19850# vss vss nfet$243
Xnfet$236_0 m1_n10452_25858# m1_n10452_25858# m1_n7186_25858# m1_n7186_25858# m1_n6629_25502#
+ vss nfet$236
Xnfet$215_5 m1_10458_17836# m1_11738_16080# m1_11271_18030# vss nfet$215
Xpfet$214_7 vdd m1_28003_18030# vdd m1_26676_16080# pfet$214
Xpfet$207_6 vdd vdd m1_31535_19792# m1_14422_22513# pfet$207
Xpfet$197_94 vdd vdd m1_22624_17518# m1_22034_17714# pfet$197
Xpfet$197_83 vdd m1_16538_15778# m1_15921_16080# m1_14641_17836# pfet$197
Xpfet$197_72 vdd m1_20721_15778# m1_20104_16080# m1_18824_17836# pfet$197
Xpfet$197_61 vdd m1_n811_16080# m1_n1278_18030# m1_n2250_17343# pfet$197
Xpfet$197_50 vdd m1_n1168_15778# m1_n1989_16202# m1_n2250_17343# pfet$197
Xpfet$205_3 vdd m1_n646_24542# vdd m1_326_24346# pfet$205
Xnfet$213_2 m1_9288_21786# m1_9288_21786# m1_9645_21447# m1_9645_21447# m1_10509_21586#
+ vss nfet$213
Xnfet$220_3 m1_n7513_20152# vss m1_326_24346# vss nfet$220
Xpfet$202_15 vdd vdd m1_22205_20152# m1_17697_15478# pfet$202
Xpfet$197_105 vdd vdd m1_14258_17518# m1_13668_17714# pfet$197
Xpfet$210_1 vdd vdd m1_34093_22102# m1_34843_21786# pfet$210
Xnfet$215_74 m1_14482_17343# vss m1_14641_17836# vss nfet$215
Xnfet$215_63 m1_13668_17714# vss m1_14258_17518# vss nfet$215
Xnfet$215_52 m1_23007_17836# m1_24287_16080# m1_23820_18030# vss nfet$215
Xnfet$215_30 sd6 vss m1_5148_15478# vss nfet$215
Xnfet$215_41 m1_n2091_17836# m1_n1168_15778# m1_n1989_16202# vss nfet$215
Xpfet$203_0 vdd vdd m1_n7401_15478# sd9 pfet$203
Xpfet$199_29 vdd vdd vdd m1_23924_19850# m1_25722_20152# m1_25722_20152# pfet$199
Xpfet$199_18 vdd vdd vdd m1_27441_19850# m1_29239_20152# m1_29239_20152# pfet$199
Xnfet$238_4 m1_2590_19404# m1_2590_19404# vss vss m1_n2445_21430# vss nfet$238
Xnfet$212_75 m1_28371_23922# vss m1_28991_24224# vss nfet$212
Xnfet$212_64 m1_19644_25858# vss m1_19781_25662# vss nfet$212
Xnfet$212_53 m1_23827_25858# m1_24451_25662# m1_24188_23922# vss nfet$212
Xnfet$212_42 m1_15943_25858# vss m1_16085_25662# vss nfet$212
Xnfet$212_31 m1_15943_25858# vss m1_18339_24542# vss nfet$212
Xnfet$217_9 m1_25747_17714# vss m1_27003_19550# vss nfet$217
Xnfet$212_20 pd3 vss m1_5771_21786# vss nfet$212
Xnfet$229_0 m1_34093_22102# vss fout vss nfet$229
Xnfet$243_2 m1_n8145_21908# vss m1_n8283_20611# vss nfet$243
Xnfet$236_1 m1_n6111_25858# m1_n6111_25858# vss vss m1_n6629_25502# vss nfet$236
Xpfet$196_19 vdd vdd m1_7095_25858# m1_4005_21786# pfet$196
Xnfet$215_6 m1_6116_17343# vss m1_6275_17836# vss nfet$215
Xpfet$207_7 vdd vdd m1_31535_22102# m1_354_22513# pfet$207
Xpfet$197_95 vdd vdd m1_21564_17714# m1_22034_17714# pfet$197
Xpfet$197_84 vdd vdd m1_17381_17714# m1_17851_17714# pfet$197
Xpfet$197_73 vdd vdd m1_16538_15778# m1_13668_17714# pfet$197
Xpfet$197_62 vdd vdd m1_23007_17836# m1_22848_17343# pfet$197
Xpfet$197_40 vdd m1_10560_16202# m1_10075_17518# m1_10458_17836# pfet$197
Xpfet$197_51 vdd vdd m1_n1168_15778# m1_n811_16080# pfet$197
Xnfet$213_3 m1_9418_21590# m1_9418_21590# m1_9645_21447# m1_9645_21447# m1_9877_21586#
+ vss nfet$213
Xnfet$220_4 m1_n789_25858# vss m1_1607_24542# vss nfet$220
Xpfet$205_4 vdd vdd m1_32675_25947# m1_33790_24346# pfet$205
Xpfet$197_106 vdd vdd m1_14482_17343# m1_17381_17714# pfet$197
Xpfet$202_16 vdd vdd m1_19969_19550# m1_17381_17714# pfet$202
Xnfet$211_0 m1_4509_24346# m1_4509_24346# vss vss m1_3991_24542# vss nfet$211
Xpfet$210_2 vdd vdd m1_30256_22102# m1_7388_22513# pfet$210
Xpfet$203_1 vdd vdd m1_21880_15478# sd2 pfet$203
Xnfet$215_31 m1_1933_17343# m1_3989_15778# m1_3372_16080# vss nfet$215
Xnfet$215_20 m1_1119_17714# vss m1_1709_17518# vss nfet$215
Xnfet$215_42 m1_n811_16080# vss m1_n1168_15778# vss nfet$215
Xnfet$215_75 sd3 vss m1_17697_15478# vss nfet$215
Xnfet$215_64 m1_13668_17714# vss m1_13198_17714# vss nfet$215
Xnfet$215_53 m1_22848_17343# vss m1_23007_17836# vss nfet$215
Xpfet$199_19 vdd m1_n3822_20130# m1_n3822_20130# m1_27441_19850# m1_27003_19550# m1_27003_19550#
+ pfet$199
Xnfet$238_5 m1_6107_19404# m1_6107_19404# m1_n5227_21418# m1_n5227_21418# m1_n2445_21430#
+ vss nfet$238
Xnfet$212_76 m1_28492_25858# vss m1_28634_25662# vss nfet$212
Xnfet$212_65 m1_28492_25858# vss m1_25107_21786# vss nfet$212
Xnfet$212_54 m1_24309_25858# vss m1_24451_25662# vss nfet$212
Xnfet$212_43 m1_15461_25858# vss m1_15598_25662# vss nfet$212
Xnfet$212_32 m1_15461_25858# m1_17546_25658# m1_18339_24542# vss nfet$212
Xnfet$212_21 m1_11278_25858# m1_11902_25662# m1_11639_23922# vss nfet$212
Xnfet$212_10 m1_7577_25858# vss m1_9973_24542# vss nfet$212
Xnfet$243_3 m1_n8283_19850# m1_n8283_20611# vss vss nfet$243
Xnfet$215_7 m1_9485_17714# vss m1_10075_17518# vss nfet$215
Xnfet$241_0 m1_n10933_25858# m1_n8848_25658# m1_n8055_24542# vss nfet$241
Xpfet$197_96 vdd vdd m1_18665_17343# m1_21564_17714# pfet$197
Xpfet$197_85 vdd m1_18926_16202# m1_18441_17518# m1_18824_17836# pfet$197
Xpfet$197_74 vdd vdd m1_14641_17836# m1_14482_17343# pfet$197
Xpfet$197_63 vdd m1_23930_15778# m1_23109_16202# m1_22848_17343# pfet$197
Xpfet$197_30 vdd vdd m1_1933_17343# m1_4832_17714# pfet$197
Xpfet$197_41 vdd vdd m1_10075_17518# m1_9485_17714# pfet$197
Xpfet$197_52 vdd m1_n3064_17714# vdd m1_n1989_16202# pfet$197
Xpfet$226_0 vdd vdd m1_n5227_20152# m1_n2543_20130# pfet$226
Xnfet$213_4 m1_5901_21590# m1_5901_21590# m1_7388_22513# m1_7388_22513# m1_6360_21586#
+ vss nfet$213
Xnfet$220_5 m1_n789_25858# vss m1_488_21786# vss nfet$220
Xpfet$205_5 vdd m1_32675_25947# vdd m1_34278_25658# pfet$205
Xnfet$220_10 m1_32675_25947# vss m1_35071_24542# vss nfet$220
Xpfet$202_17 vdd vdd m1_25722_20152# m1_21880_15478# pfet$202
Xpfet$197_107 vdd m1_15921_16080# m1_15454_18030# m1_14482_17343# pfet$197
Xpfet$203_2 vdd vdd m1_26063_15478# sd1 pfet$203
Xpfet$210_3 vdd m1_31535_22102# vdd m1_3871_22513# pfet$210
Xnfet$211_1 m1_3893_24224# m1_3893_24224# m1_3537_24542# m1_3537_24542# m1_3991_24542#
+ vss nfet$211
Xnfet$215_76 m1_14482_17343# m1_16538_15778# m1_15921_16080# vss nfet$215
Xnfet$215_65 m1_14482_17343# m1_14743_16202# m1_14258_17518# vss nfet$215
Xnfet$231_20 m1_22493_16080# m1_22493_16080# m1_22034_17714# m1_22034_17714# m1_22591_16398#
+ vss nfet$231
Xnfet$215_54 m1_22848_17343# m1_23109_16202# m1_22624_17518# vss nfet$215
Xnfet$215_32 m1_2092_17836# m1_3015_15778# m1_2194_16202# vss nfet$215
Xnfet$215_21 m1_1933_17343# m1_2194_16202# m1_1709_17518# vss nfet$215
Xnfet$215_10 m1_11738_16080# vss m1_11381_15778# vss nfet$215
Xnfet$215_43 sd8 vss m1_n3218_15478# vss nfet$215
Xnfet$238_6 m1_n5764_21786# m1_n5764_21786# vss vss m1_n6282_21430# vss nfet$238
Xnfet$212_77 m1_28010_25858# vss m1_28147_25662# vss nfet$212
Xnfet$212_66 m1_28010_25858# m1_30095_25658# m1_30888_24542# vss nfet$212
Xnfet$212_55 m1_23827_25858# vss m1_23964_25662# vss nfet$212
Xnfet$212_44 m1_15822_23922# vss m1_16442_24224# vss nfet$212
Xnfet$212_33 m1_11760_25858# vss m1_14156_24542# vss nfet$212
Xnfet$212_22 m1_11760_25858# vss m1_11902_25662# vss nfet$212
Xnfet$212_11 m1_7522_21786# vss m1_11278_25858# vss nfet$212
Xnfet$215_8 m1_7555_16080# vss m1_7198_15778# vss nfet$215
Xnfet$234_0 m1_n6274_17836# m1_n4994_16080# m1_n5461_18030# vss nfet$234
Xnfet$241_1 m1_n10796_25662# m1_n10572_23922# m1_n10308_24542# vss nfet$241
Xpfet$197_20 vdd vdd m1_1119_17714# m1_1578_16080# pfet$197
Xpfet$226_1 vdd m1_n4485_20152# vdd m1_n3206_20274# pfet$226
Xpfet$219_0 vdd vdd m1_n7320_25516# m1_n7186_25858# pfet$219
Xpfet$197_97 vdd vdd m1_22493_16080# m1_n7513_20152# pfet$197
Xpfet$197_86 vdd m1_19637_18030# vdd m1_18310_16080# pfet$197
Xpfet$197_75 vdd vdd m1_17697_15478# sd3 pfet$197
Xpfet$197_64 vdd vdd m1_23930_15778# m1_24287_16080# pfet$197
Xnfet$220_6 m1_n910_23922# vss m1_n290_24224# vss nfet$220
Xpfet$197_31 vdd m1_3372_16080# m1_2905_18030# m1_1933_17343# pfet$197
Xpfet$197_42 vdd m1_11271_18030# vdd m1_9944_16080# pfet$197
Xpfet$197_53 vdd vdd m1_n3218_15478# sd8 pfet$197
Xnfet$213_5 m1_2254_21786# m1_2254_21786# m1_3871_22513# m1_3871_22513# m1_3475_21586#
+ vss nfet$213
Xpfet$205_6 vdd vdd m1_32818_24542# m1_33174_24224# pfet$205
Xnfet$220_11 m1_32554_23922# vss m1_33174_24224# vss nfet$220
Xpfet$210_4 vdd m1_30256_22102# vdd m1_9645_21447# pfet$210
Xpfet$197_108 vdd vdd m1_15454_18030# m1_15564_15778# pfet$197
Xnfet$211_2 m1_4997_25658# m1_4997_25658# vss vss m1_5456_25502# vss nfet$211
Xnfet$215_77 sd4 vss m1_13514_15478# vss nfet$215
Xnfet$215_66 m1_n7513_20152# vss m1_14127_16080# vss nfet$215
Xnfet$231_21 m1_14127_16080# m1_14127_16080# vss vss m1_15690_17358# vss nfet$231
Xnfet$215_55 m1_22034_17714# vss m1_24904_15778# vss nfet$215
Xnfet$215_44 m1_n2091_17836# m1_n811_16080# m1_n1278_18030# vss nfet$215
Xnfet$215_33 sd7 vss m1_965_15478# vss nfet$215
Xnfet$231_10 m1_1578_16080# m1_1578_16080# m1_1119_17714# m1_1119_17714# m1_1676_16398#
+ vss nfet$231
Xnfet$215_22 m1_6116_17343# m1_6377_16202# m1_5892_17518# vss nfet$215
Xnfet$215_11 m1_10299_17343# m1_12355_15778# m1_11738_16080# vss nfet$215
Xpfet$201_0 vdd vdd m1_n6274_17836# m1_n6433_17343# pfet$201
Xnfet$238_7 m1_n3822_21786# m1_n3822_21786# m1_n4485_21904# m1_n4485_21904# m1_n3724_21430#
+ vss nfet$238
Xnfet$212_12 m1_7577_25858# vss m1_7522_21786# vss nfet$212
Xnfet$212_78 m1_28010_25858# m1_28634_25662# m1_28371_23922# vss nfet$212
Xnfet$212_67 m1_28492_25858# vss m1_30888_24542# vss nfet$212
Xnfet$212_56 m1_19781_25662# m1_20625_24224# m1_21729_25658# vss nfet$212
Xnfet$212_45 m1_15461_25858# m1_16085_25662# m1_15822_23922# vss nfet$212
Xnfet$212_34 m1_11278_25858# m1_13363_25658# m1_14156_24542# vss nfet$212
Xnfet$212_23 m1_11278_25858# vss m1_11415_25662# vss nfet$212
Xpfet$199_0 vdd m1_2590_19404# m1_2590_19404# m1_3458_19550# m1_n3534_17714# m1_n3534_17714#
+ pfet$199
Xnfet$215_9 sd5 vss m1_9331_15478# vss nfet$215
Xnfet$234_1 m1_n6433_17343# m1_n4377_15778# m1_n4994_16080# vss nfet$234
Xnfet$241_2 m1_n10933_25858# m1_n10309_25662# m1_n10572_23922# vss nfet$241
Xnfet$227_0 m1_31535_22102# m1_32818_21586# vss vss nfet$227
Xpfet$226_2 vdd m1_n5227_20152# vdd m1_n1927_20274# pfet$226
Xpfet$219_1 vdd vdd m1_n6111_25858# m1_n6856_24542# pfet$219
Xnfet$220_7 m1_25107_21786# vss m1_32193_25858# vss nfet$220
Xpfet$197_98 vdd m1_20104_16080# m1_19637_18030# m1_18665_17343# pfet$197
Xpfet$197_87 vdd vdd m1_18310_16080# m1_n7513_20152# pfet$197
Xpfet$197_76 vdd m1_17851_17714# vdd m1_18926_16202# pfet$197
Xpfet$197_65 vdd m1_24904_15778# m1_24287_16080# m1_23007_17836# pfet$197
Xpfet$197_21 vdd vdd m1_965_15478# sd7 pfet$197
Xpfet$197_10 vdd m1_8172_15778# m1_7555_16080# m1_6275_17836# pfet$197
Xpfet$197_32 vdd vdd m1_2905_18030# m1_3015_15778# pfet$197
Xpfet$197_43 vdd vdd m1_11271_18030# m1_11381_15778# pfet$197
Xpfet$197_54 vdd vdd m1_n1278_18030# m1_n1168_15778# pfet$197
Xnfet$213_6 m1_2384_21590# m1_2384_21590# m1_3871_22513# m1_3871_22513# m1_2843_21586#
+ vss nfet$213
Xpfet$205_7 vdd m1_32818_24542# vdd m1_33790_24346# pfet$205
Xnfet$220_12 m1_32675_25947# vss m1_28624_21786# vss nfet$220
Xpfet$197_109 vdd vdd m1_10299_17343# m1_13198_17714# pfet$197
Xnfet$211_3 m1_4509_24346# m1_4509_24346# m1_3394_25858# m1_3394_25858# m1_5456_25502#
+ vss nfet$211
Xnfet$215_78 m1_14641_17836# m1_15564_15778# m1_14743_16202# vss nfet$215
Xnfet$231_22 m1_15564_15778# m1_15564_15778# m1_15454_18030# m1_15454_18030# m1_15690_17358#
+ vss nfet$231
Xnfet$215_67 m1_17381_17714# vss m1_14482_17343# vss nfet$215
Xnfet$215_56 m1_24287_16080# vss m1_23930_15778# vss nfet$215
Xnfet$215_45 m1_n3064_17714# vss m1_n194_15778# vss nfet$215
Xnfet$215_34 m1_n2250_17343# vss m1_n2091_17836# vss nfet$215
Xnfet$215_23 m1_5302_17714# vss m1_4832_17714# vss nfet$215
Xnfet$215_12 m1_9485_17714# vss m1_12355_15778# vss nfet$215
Xnfet$231_11 m1_6377_16202# m1_6377_16202# vss vss m1_5859_16398# vss nfet$231
Xpfet$201_1 vdd vdd m1_n4377_15778# m1_n7247_17714# pfet$201
Xnfet$238_8 m1_9624_19404# m1_9624_19404# vss vss m1_n3724_21430# vss nfet$238
Xnfet$212_79 pd7 vss m1_19839_21786# vss nfet$212
Xnfet$212_68 m1_n7513_20152# vss m1_29607_24346# vss nfet$212
Xnfet$212_57 m1_20126_25858# vss m1_20268_25662# vss nfet$212
Xnfet$212_46 m1_20126_25858# vss m1_18073_21786# vss nfet$212
Xnfet$212_35 m1_15598_25662# m1_15822_23922# m1_16086_24542# vss nfet$212
Xnfet$212_24 m1_7095_25858# m1_7719_25662# m1_7456_23922# vss nfet$212
Xnfet$212_13 m1_11415_25662# m1_11639_23922# m1_11903_24542# vss nfet$212
Xpfet$199_1 vdd vdd vdd m1_2822_19850# m1_4620_20152# m1_4620_20152# pfet$199
Xnfet$234_2 m1_n6274_17836# m1_n5351_15778# m1_n6172_16202# vss nfet$234
Xpfet$226_3 vdd m1_n6839_20152# vdd m1_n927_19404# pfet$226
Xnfet$241_3 m1_n10796_25662# m1_n9952_24224# m1_n8848_25658# vss nfet$241
Xpfet$197_99 vdd m1_23109_16202# m1_22624_17518# m1_23007_17836# pfet$197
Xpfet$197_88 vdd vdd m1_18441_17518# m1_17851_17714# pfet$197
Xpfet$197_77 vdd vdd m1_17851_17714# m1_18310_16080# pfet$197
Xpfet$197_66 vdd vdd m1_24904_15778# m1_22034_17714# pfet$197
Xpfet$197_22 vdd vdd m1_3015_15778# m1_3372_16080# pfet$197
Xpfet$197_11 vdd vdd m1_9485_17714# m1_9944_16080# pfet$197
Xpfet$197_33 vdd vdd m1_5892_17518# m1_5302_17714# pfet$197
Xpfet$197_44 vdd vdd m1_649_17714# m1_1119_17714# pfet$197
Xpfet$197_55 vdd vdd m1_n2474_17518# m1_n3064_17714# pfet$197
Xnfet$220_8 m1_32193_25858# vss m1_32330_25662# vss nfet$220
Xnfet$213_7 m1_5771_21786# m1_5771_21786# m1_7388_22513# m1_7388_22513# m1_6992_21586#
+ vss nfet$213
Xnfet$220_13 m1_32675_25947# vss m1_32817_25662# vss nfet$220
Xpfet$224_0 vdd vdd vdd m1_n8047_19550# m1_n7513_20152# m1_n7513_20152# pfet$224
Xnfet$211_4 m1_12259_24224# m1_12259_24224# m1_11903_24542# m1_11903_24542# m1_12357_24542#
+ vss nfet$211
Xpfet$196_110 vdd m1_11903_24542# vdd m1_12875_24346# pfet$196
Xnfet$215_79 m1_15921_16080# vss m1_15564_15778# vss nfet$215
Xnfet$231_23 m1_18926_16202# m1_18926_16202# vss vss m1_18408_16398# vss nfet$231
Xnfet$215_68 m1_18665_17343# m1_18926_16202# m1_18441_17518# vss nfet$215
Xnfet$215_57 m1_22848_17343# m1_24904_15778# m1_24287_16080# vss nfet$215
Xnfet$215_46 m1_22034_17714# vss m1_21564_17714# vss nfet$215
Xnfet$215_24 m1_4832_17714# vss m1_1933_17343# vss nfet$215
Xnfet$215_13 m1_10458_17836# m1_11381_15778# m1_10560_16202# vss nfet$215
Xnfet$215_35 m1_n7513_20152# vss m1_5761_16080# vss nfet$215
Xnfet$231_12 m1_n1168_15778# m1_n1168_15778# m1_n1278_18030# m1_n1278_18030# m1_n1042_17358#
+ vss nfet$231
Xpfet$201_2 vdd vdd m1_n5351_15778# m1_n4994_16080# pfet$201
Xnfet$238_9 m1_n6380_21786# m1_n6380_21786# m1_n6839_21786# m1_n6839_21786# m1_n6282_21430#
+ vss nfet$238
Xnfet$212_69 m1_24309_25858# vss m1_26705_24542# vss nfet$212
Xnfet$212_58 m1_20005_23922# vss m1_20625_24224# vss nfet$212
Xnfet$212_47 m1_23964_25662# m1_24188_23922# m1_24452_24542# vss nfet$212
Xnfet$212_36 m1_11760_25858# vss m1_11039_21786# vss nfet$212
Xnfet$212_25 m1_7232_25662# m1_8076_24224# m1_9180_25658# vss nfet$212
Xnfet$212_14 m1_n7513_20152# vss m1_8692_24346# vss nfet$212
Xpfet$199_2 vdd m1_2590_19404# m1_2590_19404# m1_2822_19850# m1_2384_19550# m1_2384_19550#
+ pfet$199
Xnfet$234_3 m1_n6433_17343# m1_n6172_16202# m1_n6657_17518# vss nfet$234
Xnfet$241_4 m1_n4623_25487# m1_n2567_23922# m1_n3184_24224# vss nfet$241
Xpfet$197_89 vdd vdd m1_22848_17343# m1_25747_17714# pfet$197
Xpfet$197_78 vdd vdd m1_13514_15478# sd4 pfet$197
Xpfet$197_67 vdd m1_22034_17714# vdd m1_23109_16202# pfet$197
Xpfet$197_12 vdd m1_3989_15778# m1_3372_16080# m1_2092_17836# pfet$197
Xpfet$197_23 vdd m1_5302_17714# vdd m1_6377_16202# pfet$197
Xpfet$197_34 vdd vdd m1_5761_16080# m1_n7513_20152# pfet$197
Xpfet$197_45 vdd vdd m1_9944_16080# m1_n7513_20152# pfet$197
Xpfet$226_4 vdd vdd m1_n6839_20152# m1_n6973_21481# pfet$226
Xpfet$197_56 vdd m1_n1278_18030# vdd m1_n2605_16080# pfet$197
Xnfet$220_9 m1_n7513_20152# vss m1_33790_24346# vss nfet$220
Xnfet$213_8 m1_23486_21590# m1_23486_21590# m1_24973_22513# m1_24973_22513# m1_23945_21586#
+ vss nfet$213
Xnfet$232_0 m1_4620_20152# m1_4620_20152# m1_2590_19404# m1_2590_19404# m1_3454_20470#
+ vss nfet$232
Xpfet$224_1 vdd m1_n8283_19850# m1_n8283_19850# m1_n8047_19550# m1_n8283_20611# m1_n8283_20611#
+ pfet$224
Xpfet$217_0 vdd vdd vdd m1_n6624_23622# m1_n7082_23622# m1_n7082_23622# pfet$217
Xnfet$211_5 m1_8692_24346# m1_8692_24346# vss vss m1_8174_24542# vss nfet$211
Xpfet$196_100 vdd vdd m1_29607_24346# m1_n7513_20152# pfet$196
Xnfet$215_58 m1_23007_17836# m1_23930_15778# m1_23109_16202# vss nfet$215
Xnfet$215_47 m1_22034_17714# vss m1_22624_17518# vss nfet$215
Xnfet$215_25 m1_2092_17836# m1_3372_16080# m1_2905_18030# vss nfet$215
Xnfet$215_14 m1_6116_17343# m1_8172_15778# m1_7555_16080# vss nfet$215
Xnfet$215_36 m1_n3064_17714# vss m1_n2474_17518# vss nfet$215
Xnfet$231_24 m1_18310_16080# m1_18310_16080# m1_17851_17714# m1_17851_17714# m1_18408_16398#
+ vss nfet$231
Xnfet$215_69 m1_17851_17714# vss m1_17381_17714# vss nfet$215
Xnfet$231_13 m1_n2605_16080# m1_n2605_16080# vss vss m1_n1042_17358# vss nfet$231
Xpfet$201_3 vdd vdd m1_n6657_17518# m1_n7247_17714# pfet$201
Xnfet$212_59 m1_19644_25858# m1_20268_25662# m1_20005_23922# vss nfet$212
Xnfet$212_48 m1_18073_21786# vss m1_23827_25858# vss nfet$212
Xnfet$212_37 m1_11039_21786# vss m1_15461_25858# vss nfet$212
Xnfet$212_26 m1_7095_25858# m1_9180_25658# m1_9973_24542# vss nfet$212
Xnfet$212_15 m1_7232_25662# m1_7456_23922# m1_7720_24542# vss nfet$212
Xpfet$200_10 vdd vdd m1_23486_21590# m1_23356_21786# pfet$200
Xpfet$199_3 vdd vdd vdd m1_3458_19550# m1_n3218_15478# m1_n3218_15478# pfet$199
Xnfet$234_4 m1_27031_17343# m1_27292_16202# m1_26807_17518# vss nfet$234
Xnfet$241_5 m1_n4464_25980# m1_n3541_23922# m1_n4362_24346# vss nfet$241
Xpfet$197_79 vdd m1_15564_15778# m1_14743_16202# m1_14482_17343# pfet$197
Xpfet$197_68 vdd vdd m1_22034_17714# m1_22493_16080# pfet$197
Xpfet$197_13 vdd vdd m1_5148_15478# sd6 pfet$197
Xpfet$197_0 vdd vdd m1_12355_15778# m1_9485_17714# pfet$197
Xpfet$197_24 vdd m1_6377_16202# m1_5892_17518# m1_6275_17836# pfet$197
Xpfet$197_35 vdd vdd m1_9015_17714# m1_9485_17714# pfet$197
Xpfet$197_46 vdd vdd m1_n2250_17343# m1_649_17714# pfet$197
Xpfet$197_57 vdd m1_n1989_16202# m1_n2474_17518# m1_n2091_17836# pfet$197
Xnfet$213_9 m1_23356_21786# m1_23356_21786# m1_24973_22513# m1_24973_22513# m1_24577_21586#
+ vss nfet$213
Xnfet$225_0 m1_21456_22513# m1_21456_22513# m1_30256_19792# m1_30256_19792# m1_30492_20470#
+ vss nfet$225
Xnfet$232_1 m1_1103_20152# m1_1103_20152# m1_n927_19404# m1_n927_19404# m1_n63_20470#
+ vss nfet$232
Xpfet$224_2 vdd m1_n8283_20611# m1_n8283_20611# m1_n8047_22344# m1_n8145_21908# m1_n8145_21908#
+ pfet$224
Xpfet$217_1 vdd m1_n6856_24542# m1_n6856_24542# m1_n6624_23622# m1_n8283_19850# m1_n8283_19850#
+ pfet$217
Xpfet$196_101 vdd vdd m1_28010_25858# m1_21590_21786# pfet$196
Xnfet$211_6 m1_8076_24224# m1_8076_24224# m1_7720_24542# m1_7720_24542# m1_8174_24542#
+ vss nfet$211
Xnfet$231_25 m1_14743_16202# m1_14743_16202# vss vss m1_14225_16398# vss nfet$231
Xnfet$215_59 m1_17851_17714# vss m1_20721_15778# vss nfet$215
Xnfet$215_48 m1_18824_17836# m1_20104_16080# m1_19637_18030# vss nfet$215
Xnfet$215_26 m1_5302_17714# vss m1_5892_17518# vss nfet$215
Xnfet$215_15 m1_5302_17714# vss m1_8172_15778# vss nfet$215
Xnfet$215_37 m1_n7513_20152# vss m1_n2605_16080# vss nfet$215
Xnfet$231_14 m1_n2605_16080# m1_n2605_16080# m1_n3064_17714# m1_n3064_17714# m1_n2507_16398#
+ vss nfet$231
Xpfet$201_4 vdd vdd m1_n6433_17343# m1_n3534_17714# pfet$201
Xnfet$212_49 m1_19781_25662# m1_20005_23922# m1_20269_24542# vss nfet$212
Xnfet$212_38 m1_n7513_20152# vss m1_12875_24346# vss nfet$212
Xnfet$212_27 m1_7577_25858# vss m1_7719_25662# vss nfet$212
Xnfet$212_16 m1_4005_21786# vss m1_7095_25858# vss nfet$212
Xpfet$200_11 vdd vdd m1_18705_21786# m1_18073_21786# pfet$200
Xpfet$199_4 vdd m1_6107_19404# m1_6107_19404# m1_6339_19850# m1_5901_19550# m1_5901_19550#
+ pfet$199
Xnfet$234_5 m1_27031_17343# m1_29087_15778# m1_28470_16080# vss nfet$234
Xnfet$241_6 m1_n4464_25980# m1_n3184_24224# m1_n3651_26174# vss nfet$241
Xpfet$197_14 vdd vdd m1_2092_17836# m1_1933_17343# pfet$197
Xpfet$197_1 vdd vdd m1_11381_15778# m1_11738_16080# pfet$197
Xpfet$197_25 vdd vdd m1_1709_17518# m1_1119_17714# pfet$197
Xpfet$197_36 vdd vdd m1_6116_17343# m1_9015_17714# pfet$197
Xpfet$197_69 vdd vdd m1_20721_15778# m1_17851_17714# pfet$197
Xpfet$197_47 vdd m1_11738_16080# m1_11271_18030# m1_10299_17343# pfet$197
Xpfet$197_58 vdd vdd m1_n3534_17714# m1_n3064_17714# pfet$197
Xnfet$225_1 m1_14422_22513# m1_14422_22513# m1_31535_19792# m1_31535_19792# m1_31771_20470#
+ vss nfet$225
Xnfet$232_2 m1_n3218_15478# m1_n3218_15478# m1_2590_19404# m1_2590_19404# m1_2822_20470#
+ vss nfet$232
Xnfet$218_0 sd9 vss m1_n7401_15478# vss nfet$218
Xpfet$224_3 vdd vdd vdd m1_n8047_22344# m1_n8283_19850# m1_n8283_19850# pfet$224
Xnfet$211_7 m1_9180_25658# m1_9180_25658# vss vss m1_9639_25502# vss nfet$211
Xpfet$196_102 vdd m1_28371_23922# m1_28635_24542# m1_28010_25858# pfet$196
Xnfet$231_26 m1_14127_16080# m1_14127_16080# m1_13668_17714# m1_13668_17714# m1_14225_16398#
+ vss nfet$231
Xnfet$215_49 m1_21564_17714# vss m1_18665_17343# vss nfet$215
Xnfet$215_27 m1_1119_17714# vss m1_3989_15778# vss nfet$215
Xnfet$215_16 m1_6275_17836# m1_7198_15778# m1_6377_16202# vss nfet$215
Xnfet$215_38 m1_n2250_17343# m1_n1989_16202# m1_n2474_17518# vss nfet$215
Xnfet$231_15 m1_n1989_16202# m1_n1989_16202# vss vss m1_n2507_16398# vss nfet$231
Xpfet$222_0 vdd vdd m1_n10796_25662# m1_n10933_25858# pfet$222
Xpfet$201_5 vdd vdd m1_n6788_16080# m1_n7513_20152# pfet$201
Xnfet$212_28 m1_3394_25858# vss m1_4005_21786# vss nfet$212
Xnfet$212_17 m1_11639_23922# vss m1_12259_24224# vss nfet$212
Xnfet$212_39 pd4 vss m1_9288_21786# vss nfet$212
Xpfet$200_12 vdd vdd m1_16452_21590# m1_16322_21786# pfet$200
Xpfet$199_5 vdd vdd vdd m1_n695_19850# m1_1103_20152# m1_1103_20152# pfet$199
Xnfet$234_6 m1_27190_17836# m1_28113_15778# m1_27292_16202# vss nfet$234
Xnfet$241_7 m1_n4623_25487# m1_n4362_24346# m1_n4847_25662# vss nfet$241
Xpfet$197_15 vdd vdd m1_5302_17714# m1_5761_16080# pfet$197
Xpfet$197_2 vdd m1_12355_15778# m1_11738_16080# m1_10458_17836# pfet$197
Xpfet$197_26 vdd vdd m1_4832_17714# m1_5302_17714# pfet$197
Xpfet$197_37 vdd m1_7555_16080# m1_7088_18030# m1_6116_17343# pfet$197
Xpfet$197_48 vdd vdd m1_n3064_17714# m1_n2605_16080# pfet$197
Xpfet$197_59 vdd vdd m1_n2605_16080# m1_n7513_20152# pfet$197
Xnfet$218_1 sd2 vss m1_21880_15478# vss nfet$218
Xnfet$225_2 m1_17939_22513# m1_17939_22513# vss vss m1_31771_20470# vss nfet$225
Xnfet$232_3 m1_8137_20152# m1_8137_20152# m1_6107_19404# m1_6107_19404# m1_6971_20470#
+ vss nfet$232
Xpfet$222_10 vdd vdd m1_n10933_25858# fin pfet$222
Xnfet$211_8 m1_8692_24346# m1_8692_24346# m1_7577_25858# m1_7577_25858# m1_9639_25502#
+ vss nfet$211
Xpfet$196_103 vdd vdd m1_28635_24542# m1_28991_24224# pfet$196
Xnfet$230_0 fout vss m1_35837_22102# vss nfet$230
Xnfet$231_27 m1_18310_16080# m1_18310_16080# vss vss m1_19873_17358# vss nfet$231
Xnfet$231_16 m1_19747_15778# m1_19747_15778# m1_19637_18030# m1_19637_18030# m1_19873_17358#
+ vss nfet$231
Xnfet$215_28 m1_1933_17343# vss m1_2092_17836# vss nfet$215
Xnfet$215_17 m1_649_17714# vss m1_n2250_17343# vss nfet$215
Xnfet$215_39 m1_n3064_17714# vss m1_n3534_17714# vss nfet$215
Xpfet$222_1 vdd vdd m1_n10309_25662# m1_n10452_25858# pfet$222
Xpfet$215_0 vdd m1_n4377_15778# m1_n4994_16080# m1_n6274_17836# pfet$215
Xpfet$201_6 vdd vdd m1_n7383_17599# m1_n7247_17714# pfet$201
Xnfet$212_29 m1_15943_25858# vss m1_14556_21786# vss nfet$212
Xnfet$212_18 m1_7095_25858# vss m1_7232_25662# vss nfet$212
Xpfet$200_13 vdd vdd m1_15188_21786# m1_14556_21786# pfet$200
Xpfet$199_6 vdd vdd vdd m1_6339_19850# m1_8137_20152# m1_8137_20152# pfet$199
Xnfet$234_7 m1_27190_17836# m1_28470_16080# m1_28003_18030# vss nfet$234
Xpfet$197_16 vdd vdd m1_3989_15778# m1_1119_17714# pfet$197
Xpfet$197_3 vdd m1_11381_15778# m1_10560_16202# m1_10299_17343# pfet$197
Xpfet$197_27 vdd m1_2194_16202# m1_1709_17518# m1_2092_17836# pfet$197
Xpfet$197_38 vdd vdd m1_7088_18030# m1_7198_15778# pfet$197
Xpfet$197_49 vdd m1_n194_15778# m1_n811_16080# m1_n2091_17836# pfet$197
Xnfet$218_2 sd1 vss m1_26063_15478# vss nfet$218
Xnfet$225_3 m1_24973_22513# m1_24973_22513# vss vss m1_30492_20470# vss nfet$225
Xnfet$232_4 m1_965_15478# m1_965_15478# m1_6107_19404# m1_6107_19404# m1_6339_20470#
+ vss nfet$232
Xpfet$222_11 vdd vdd m1_n9336_24346# vss pfet$222
Xnfet$211_9 m1_17058_24346# m1_17058_24346# vss vss m1_16540_24542# vss nfet$211
Xpfet$196_104 vdd m1_25912_25658# m1_26705_24542# m1_23964_25662# pfet$196
Xnfet$230_1 define m1_35837_22102# vss vss nfet$230
Xnfet$231_17 m1_22493_16080# m1_22493_16080# vss vss m1_24056_17358# vss nfet$231
Xnfet$215_29 m1_3372_16080# vss m1_3015_15778# vss nfet$215
Xnfet$215_18 m1_1119_17714# vss m1_649_17714# vss nfet$215
Xnfet$223_0 m1_n290_24224# m1_n290_24224# m1_n646_24542# m1_n646_24542# m1_n192_24542#
+ vss nfet$223
Xpfet$215_1 vdd m1_n5351_15778# m1_n6172_16202# m1_n6433_17343# pfet$215
Xpfet$222_2 vdd vdd m1_n9952_24224# m1_n10572_23922# pfet$222
Xpfet$208_0 vdd m1_n647_25662# m1_n910_23922# m1_n1134_25662# pfet$208
Xpfet$201_7 vdd vdd m1_27190_17836# m1_27031_17343# pfet$201
Xnfet$212_19 m1_7456_23922# vss m1_8076_24224# vss nfet$212
Xpfet$200_14 vdd vdd m1_19969_21590# m1_19839_21786# pfet$200
Xpfet$199_7 vdd vdd vdd m1_6975_19550# m1_965_15478# m1_965_15478# pfet$199
Xpfet$197_17 vdd vdd m1_n2091_17836# m1_n2250_17343# pfet$197
Xpfet$197_4 vdd m1_9485_17714# vdd m1_10560_16202# pfet$197
Xpfet$197_28 vdd m1_2905_18030# vdd m1_1578_16080# pfet$197
Xpfet$197_39 vdd m1_7088_18030# vdd m1_5761_16080# pfet$197
Xnfet$225_4 m1_32818_20470# m1_32818_20470# vss vss m1_34329_20470# vss nfet$225
Xnfet$232_5 m1_5148_15478# m1_5148_15478# m1_9624_19404# m1_9624_19404# m1_9856_20470#
+ vss nfet$232
Xpfet$222_12 vdd vdd m1_n7082_23622# m1_n8625_26174# pfet$222
Xpfet$196_105 vdd vdd m1_30888_24542# m1_28492_25858# pfet$196
Xnfet$223_1 m1_814_25658# m1_814_25658# vss vss m1_1273_25502# vss nfet$223
Xnfet$215_19 m1_n7513_20152# vss m1_1578_16080# vss nfet$215
Xnfet$216_0 m1_n1263_21786# vss m1_n1133_21590# vss nfet$216
Xnfet$231_18 m1_23930_15778# m1_23930_15778# m1_23820_18030# m1_23820_18030# m1_24056_17358#
+ vss nfet$231
Xpfet$215_2 vdd m1_n4994_16080# m1_n5461_18030# m1_n6433_17343# pfet$215
Xpfet$222_3 vdd vdd m1_n4978_24224# vss pfet$222
Xpfet$208_1 vdd m1_n910_23922# m1_n646_24542# m1_n1271_25858# pfet$208
Xpfet$201_8 vdd vdd m1_28113_15778# m1_28470_16080# pfet$201
Xpfet$220_0 vdd vdd m1_n8625_26174# m1_n9336_24346# pfet$220
Xpfet$200_15 vdd vdd m1_27003_21590# m1_26873_21786# pfet$200
Xpfet$199_8 vdd m1_9624_19404# m1_9624_19404# m1_10492_19550# m1_4832_17714# m1_4832_17714#
+ pfet$199
Xpfet$197_18 vdd m1_1119_17714# vdd m1_2194_16202# pfet$197
Xpfet$197_5 vdd m1_7198_15778# m1_6377_16202# m1_6116_17343# pfet$197
Xpfet$197_29 vdd vdd m1_1578_16080# m1_n7513_20152# pfet$197
Xnfet$246_0 m1_n4485_20152# m1_n6380_21786# vss vss nfet$246
Xnfet$225_5 m1_32818_21586# m1_32818_21586# m1_34093_19792# m1_34093_19792# m1_34329_20470#
+ vss nfet$225
Xnfet$232_6 m1_11654_20152# m1_11654_20152# m1_9624_19404# m1_9624_19404# m1_10488_20470#
+ vss nfet$232
Xpfet$222_13 vdd vdd m1_n8055_24542# m1_n8625_26174# pfet$222
Xpfet$196_106 vdd vdd m1_25107_21786# m1_28492_25858# pfet$196
Xnfet$223_2 m1_326_24346# m1_326_24346# m1_n789_25858# m1_n789_25858# m1_1273_25502#
+ vss nfet$223
Xnfet$231_19 m1_23109_16202# m1_23109_16202# vss vss m1_22591_16398# vss nfet$231
Xpfet$215_3 vdd m1_n6172_16202# m1_n6657_17518# m1_n6274_17836# pfet$215
Xpfet$222_4 vdd vdd m1_n5571_25662# m1_n10452_25858# pfet$222
Xnfet$216_1 m1_11039_21786# vss m1_11671_21786# vss nfet$216
Xpfet$208_2 vdd m1_n290_24224# m1_814_25658# m1_n1271_25858# pfet$208
Xpfet$201_9 vdd vdd m1_29087_15778# m1_26217_17714# pfet$201
Xpfet$213_0 vdd m1_32818_20470# m1_32818_20470# m1_33050_19550# m1_30256_19792# m1_30256_19792#
+ pfet$213
Xpfet$220_1 vdd m1_n8625_26174# vdd m1_n8848_25658# pfet$220
Xpfet$200_16 vdd vdd m1_29256_21786# m1_28624_21786# pfet$200
Xpfet$199_9 vdd m1_9624_19404# m1_9624_19404# m1_9856_19850# m1_9418_19550# m1_9418_19550#
+ pfet$199
Xpfet$197_19 vdd m1_3015_15778# m1_2194_16202# m1_1933_17343# pfet$197
Xpfet$197_6 vdd vdd m1_7198_15778# m1_7555_16080# pfet$197
Xnfet$246_1 m1_n5227_20152# vss m1_n6380_21786# vss nfet$246
Xnfet$239_0 m1_n8625_26174# vss m1_n8055_24542# vss nfet$239
Xnfet$225_6 m1_354_22513# m1_354_22513# m1_31535_22102# m1_31535_22102# m1_31771_21430#
+ vss nfet$225
Xnfet$232_7 m1_n7401_15478# m1_n7401_15478# m1_n927_19404# m1_n927_19404# m1_n695_20470#
+ vss nfet$232
Xpfet$196_107 vdd m1_24309_25858# vdd m1_25912_25658# pfet$196
Xpfet$215_4 vdd m1_28113_15778# m1_27292_16202# m1_27031_17343# pfet$215
Xnfet$223_3 m1_326_24346# m1_326_24346# vss vss m1_n192_24542# vss nfet$223
Xpfet$208_3 vdd m1_814_25658# m1_1607_24542# m1_n1134_25662# pfet$208
Xpfet$222_5 vdd vdd m1_n4847_25662# m1_n10452_25858# pfet$222
Xnfet$216_2 m1_12805_21786# vss m1_12935_21590# vss nfet$216
Xnfet$221_0 m1_n1134_25662# m1_n910_23922# m1_n646_24542# vss nfet$221
Xpfet$206_0 vdd vdd vdd m1_33050_22344# m1_31535_22102# m1_31535_22102# pfet$206
Xpfet$213_1 vdd vdd vdd m1_33050_19550# m1_31535_19792# m1_31535_19792# pfet$213
Xpfet$220_2 vdd m1_n3651_26174# vdd m1_n4978_24224# pfet$220
Xpfet$200_17 vdd vdd m1_25739_21786# m1_25107_21786# pfet$200
Xnfet$213_10 m1_19839_21786# m1_19839_21786# m1_21456_22513# m1_21456_22513# m1_21060_21586#
+ vss nfet$213
Xnfet$239_1 m1_n8625_26174# vss m1_n7082_23622# vss nfet$239
Xpfet$197_7 vdd vdd m1_6275_17836# m1_6116_17343# pfet$197
Xnfet$225_7 m1_3871_22513# m1_3871_22513# vss vss m1_31771_21430# vss nfet$225
Xnfet$232_8 m1_26063_15478# m1_26063_15478# m1_n3822_20130# m1_n3822_20130# m1_27441_20470#
+ vss nfet$232
Xpfet$198_30 vdd vdd vdd m1_17539_22402# m1_16322_21786# m1_16322_21786# pfet$198
Xpfet$196_108 vdd vdd m1_25424_24346# m1_n7513_20152# pfet$196
Xnfet$223_4 m1_33174_24224# m1_33174_24224# m1_32818_24542# m1_32818_24542# m1_33272_24542#
+ vss nfet$223
Xpfet$222_6 vdd vdd m1_n4623_25487# fin pfet$222
Xnfet$216_3 m1_9288_21786# vss m1_9418_21590# vss nfet$216
Xpfet$208_4 vdd m1_33174_24224# m1_34278_25658# m1_32193_25858# pfet$208
Xpfet$215_5 vdd m1_29087_15778# m1_28470_16080# m1_27190_17836# pfet$215
Xpfet$213_2 vdd m1_32818_21586# m1_32818_21586# m1_33050_22344# m1_30256_22102# m1_30256_22102#
+ pfet$213
Xnfet$216_10 m1_21590_21786# vss m1_22222_21786# vss nfet$216
Xnfet$214_0 m1_n3534_17714# m1_n3534_17714# vss vss m1_3454_20470# vss nfet$214
Xnfet$221_1 m1_n1271_25858# m1_n647_25662# m1_n910_23922# vss nfet$221
Xpfet$220_3 vdd vdd m1_n3651_26174# m1_n3541_23922# pfet$220
Xnfet$213_11 m1_19969_21590# m1_19969_21590# m1_21456_22513# m1_21456_22513# m1_20428_21586#
+ vss nfet$213
Xpfet$197_8 vdd vdd m1_9331_15478# sd5 pfet$197
Xnfet$239_2 vss vss m1_n9336_24346# vss nfet$239
Xnfet$224_10 m1_21590_21786# m1_21590_21786# vss vss m1_20428_21586# vss nfet$224
Xnfet$232_9 m1_29239_20152# m1_29239_20152# m1_n3822_20130# m1_n3822_20130# m1_28073_20470#
+ vss nfet$232
Xnfet$244_0 m1_n4485_21904# m1_n5764_21786# vss vss nfet$244
Xpfet$198_31 vdd vdd vdd m1_27462_22102# m1_27003_21590# m1_27003_21590# pfet$198
Xpfet$198_20 vdd vdd vdd m1_20428_22102# m1_19969_21590# m1_19969_21590# pfet$198
Xnfet$219_10 m1_26217_17714# vss m1_29087_15778# vss nfet$219
Xpfet$196_109 vdd m1_12259_24224# m1_13363_25658# m1_11278_25858# pfet$196
Xnfet$223_5 m1_33790_24346# m1_33790_24346# vss vss m1_33272_24542# vss nfet$223
Xnfet$216_4 m1_7522_21786# vss m1_8154_21786# vss nfet$216
Xpfet$208_5 vdd m1_32817_25662# m1_32554_23922# m1_32330_25662# pfet$208
Xpfet$215_6 vdd m1_28470_16080# m1_28003_18030# m1_27031_17343# pfet$215
Xpfet$222_7 vdd vdd m1_n3541_23922# m1_n3184_24224# pfet$222
Xnfet$214_1 m1_2384_19550# m1_2384_19550# vss vss m1_2822_20470# vss nfet$214
Xpfet$220_4 vdd m1_n10452_25858# vdd m1_n4362_24346# pfet$220
Xnfet$221_2 m1_n1271_25858# m1_814_25658# m1_1607_24542# vss nfet$221
Xnfet$216_11 m1_18073_21786# vss m1_18705_21786# vss nfet$216
Xnfet$232_10 m1_9331_15478# m1_9331_15478# m1_n3822_21786# m1_n3822_21786# m1_13373_20470#
+ vss nfet$232
Xpfet$211_0 vdd vdd vdd m1_36073_22344# define define pfet$211
Xnfet$213_12 m1_16322_21786# m1_16322_21786# m1_17939_22513# m1_17939_22513# m1_17543_21586#
+ vss nfet$213
Xpfet$197_9 vdd vdd m1_8172_15778# m1_5302_17714# pfet$197
Xnfet$239_3 fin vss m1_n10933_25858# vss nfet$239
Xnfet$224_11 m1_22222_21786# m1_22222_21786# vss vss m1_21060_21586# vss nfet$224
Xnfet$244_1 m1_n5227_21418# vss m1_n5764_21786# vss nfet$244
Xnfet$237_0 m1_n7082_23622# m1_n6856_24542# vss vss nfet$237
Xnfet$219_11 m1_27031_17343# vss m1_27190_17836# vss nfet$219
Xnfet$223_6 m1_33790_24346# m1_33790_24346# m1_32675_25947# m1_32675_25947# m1_34737_25502#
+ vss nfet$223
Xpfet$198_32 vdd m1_28490_22513# m1_28490_22513# m1_28090_22402# m1_28624_21786# m1_28624_21786#
+ pfet$198
Xpfet$198_21 vdd vdd vdd m1_21056_22402# m1_19839_21786# m1_19839_21786# pfet$198
Xnfet$216_5 m1_488_21786# vss m1_1120_21786# vss nfet$216
Xpfet$198_10 vdd m1_3871_22513# m1_3871_22513# m1_2843_22102# m1_4637_21786# m1_4637_21786#
+ pfet$198
Xpfet$208_6 vdd m1_34278_25658# m1_35071_24542# m1_32330_25662# pfet$208
Xpfet$215_7 vdd m1_27292_16202# m1_26807_17518# m1_27190_17836# pfet$215
Xpfet$222_8 vdd vdd m1_n2567_23922# m1_n7320_25516# pfet$222
Xnfet$221_3 m1_n1134_25662# m1_n290_24224# m1_814_25658# vss nfet$221
Xnfet$214_2 m1_5901_19550# m1_5901_19550# vss vss m1_6339_20470# vss nfet$214
Xnfet$216_12 m1_14556_21786# vss m1_15188_21786# vss nfet$216
Xnfet$232_11 m1_15171_20152# m1_15171_20152# m1_n3822_21786# m1_n3822_21786# m1_14005_20470#
+ vss nfet$232
Xpfet$220_5 vdd vdd m1_n10308_24542# m1_n9952_24224# pfet$220
Xpfet$211_1 vdd m1_35837_22102# m1_35837_22102# m1_36073_22344# fout fout pfet$211
Xpfet$204_0 vdd vdd m1_n647_25662# m1_n789_25858# pfet$204
Xnfet$213_13 m1_16452_21590# m1_16452_21590# m1_17939_22513# m1_17939_22513# m1_16911_21586#
+ vss nfet$213
Xnfet$239_4 m1_n10572_23922# vss m1_n9952_24224# vss nfet$239
Xnfet$224_12 m1_18073_21786# m1_18073_21786# vss vss m1_16911_21586# vss nfet$224
Xnfet$219_12 m1_28470_16080# vss m1_28113_15778# vss nfet$219
Xnfet$244_2 m1_n6839_21786# vss m1_n6973_21481# vss nfet$244
Xnfet$237_1 m1_n8283_19850# vss m1_n6856_24542# vss nfet$237
Xnfet$223_7 m1_34278_25658# m1_34278_25658# vss vss m1_34737_25502# vss nfet$223
Xpfet$198_33 vdd m1_28490_22513# m1_28490_22513# m1_27462_22102# m1_29256_21786# m1_29256_21786#
+ pfet$198
Xpfet$198_22 vdd m1_21456_22513# m1_21456_22513# m1_20428_22102# m1_22222_21786# m1_22222_21786#
+ pfet$198
Xpfet$198_11 vdd vdd vdd m1_2843_22102# m1_2384_21590# m1_2384_21590# pfet$198
Xpfet$208_7 vdd m1_32554_23922# m1_32818_24542# m1_32193_25858# pfet$208
Xpfet$222_9 vdd vdd m1_n4464_25980# m1_n4623_25487# pfet$222
Xnfet$216_6 m1_5771_21786# vss m1_5901_21590# vss nfet$216
Xnfet$221_4 m1_32193_25858# m1_34278_25658# m1_35071_24542# vss nfet$221
Xnfet$214_3 m1_4832_17714# m1_4832_17714# vss vss m1_10488_20470# vss nfet$214
Xnfet$216_13 m1_16322_21786# vss m1_16452_21590# vss nfet$216
Xnfet$232_12 m1_18688_20152# m1_18688_20152# m1_n1927_20274# m1_n1927_20274# m1_17522_20470#
+ vss nfet$232
Xpfet$220_6 vdd m1_n10308_24542# vdd m1_n9336_24346# pfet$220
Xnfet$212_0 m1_3394_25858# vss m1_5790_24542# vss nfet$212
Xpfet$204_1 vdd vdd m1_n1134_25662# m1_n1271_25858# pfet$204
Xnfet$213_14 m1_12805_21786# m1_12805_21786# m1_14422_22513# m1_14422_22513# m1_14026_21586#
+ vss nfet$213
Xnfet$239_5 m1_n10933_25858# vss m1_n10796_25662# vss nfet$239
Xnfet$224_13 m1_18705_21786# m1_18705_21786# vss vss m1_17543_21586# vss nfet$224
Xnfet$219_13 m1_26217_17714# vss m1_25747_17714# vss nfet$219
Xpfet$198_34 vdd vdd vdd m1_28090_22402# m1_26873_21786# m1_26873_21786# pfet$198
Xpfet$198_23 vdd vdd vdd m1_23945_22102# m1_23486_21590# m1_23486_21590# pfet$198
Xpfet$198_12 vdd vdd vdd m1_3471_22402# m1_2254_21786# m1_2254_21786# pfet$198
Xnfet$242_0 m1_n7186_25858# vss m1_n7320_25516# vss nfet$242
Xnfet$216_7 m1_4005_21786# vss m1_4637_21786# vss nfet$216
Xpfet$227_0 vdd vdd vdd m1_n5019_19550# m1_n4485_20152# m1_n4485_20152# pfet$227
Xnfet$221_5 m1_32330_25662# m1_33174_24224# m1_34278_25658# vss nfet$221
Xnfet$214_4 m1_9418_19550# m1_9418_19550# vss vss m1_9856_20470# vss nfet$214
Xnfet$216_14 m1_19839_21786# vss m1_19969_21590# vss nfet$216
Xnfet$232_13 m1_13514_15478# m1_13514_15478# m1_n1927_20274# m1_n1927_20274# m1_16890_20470#
+ vss nfet$232
Xpfet$220_7 vdd vdd m1_n10452_25858# m1_n4978_24224# pfet$220
Xnfet$212_1 m1_2912_25858# m1_4997_25658# m1_5790_24542# vss nfet$212
Xpfet$204_2 vdd vdd m1_n1271_25858# m1_n10452_25858# pfet$204
Xnfet$213_15 m1_26873_21786# m1_26873_21786# m1_28490_22513# m1_28490_22513# m1_28094_21586#
+ vss nfet$213
Xnfet$239_6 m1_n10452_25858# vss m1_n10309_25662# vss nfet$239
Xnfet$224_14 m1_15188_21786# m1_15188_21786# vss vss m1_14026_21586# vss nfet$224
Xpfet$201_10 vdd vdd m1_27031_17343# m1_n10452_25858# pfet$201
Xpfet$198_35 vdd vdd vdd m1_13394_22102# m1_12935_21590# m1_12935_21590# pfet$198
Xpfet$198_24 vdd m1_17939_22513# m1_17939_22513# m1_16911_22102# m1_18705_21786# m1_18705_21786#
+ pfet$198
Xpfet$198_13 vdd vdd vdd m1_6988_22402# m1_5771_21786# m1_5771_21786# pfet$198
Xnfet$216_8 m1_2254_21786# vss m1_2384_21590# vss nfet$216
Xnfet$235_0 m1_n5351_15778# m1_n5351_15778# m1_n5461_18030# m1_n5461_18030# m1_n5225_17358#
+ vss nfet$235
Xnfet$242_1 m1_n6856_24542# vss m1_n6111_25858# vss nfet$242
Xnfet$221_6 m1_32193_25858# m1_32817_25662# m1_32554_23922# vss nfet$221
Xnfet$216_15 m1_28624_21786# vss m1_29256_21786# vss nfet$216
Xnfet$214_5 m1_649_17714# m1_649_17714# vss vss m1_6971_20470# vss nfet$214
Xnfet$232_14 m1_22205_20152# m1_22205_20152# m1_n2543_20130# m1_n2543_20130# m1_21039_20470#
+ vss nfet$232
Xpfet$204_10 vdd vdd m1_35071_24542# m1_32675_25947# pfet$204
Xnfet$212_2 m1_n7513_20152# vss m1_4509_24346# vss nfet$212
Xpfet$204_3 vdd vdd m1_1607_24542# m1_n789_25858# pfet$204
Xpfet$196_90 vdd vdd m1_24309_25858# m1_25424_24346# pfet$196
Xnfet$213_16 m1_27003_21590# m1_27003_21590# m1_28490_22513# m1_28490_22513# m1_27462_21586#
+ vss nfet$213
Xpfet$202_0 vdd vdd m1_2384_19550# m1_n3534_17714# pfet$202
Xpfet$201_11 vdd vdd m1_26807_17518# m1_26217_17714# pfet$201
Xnfet$239_7 m1_n7320_25516# vss m1_n2567_23922# vss nfet$239
Xnfet$224_15 m1_14556_21786# m1_14556_21786# vss vss m1_13394_21586# vss nfet$224
Xpfet$198_25 vdd m1_17939_22513# m1_17939_22513# m1_17539_22402# m1_18073_21786# m1_18073_21786#
+ pfet$198
Xpfet$198_14 vdd vdd vdd m1_n46_22402# m1_n1263_21786# m1_n1263_21786# pfet$198
Xnfet$216_9 m1_23356_21786# vss m1_23486_21590# vss nfet$216
Xnfet$228_0 m1_34093_19792# vss m1_34843_21786# vss nfet$228
Xnfet$235_1 m1_n6788_16080# m1_n6788_16080# vss vss m1_n5225_17358# vss nfet$235
Xnfet$221_7 m1_32330_25662# m1_32554_23922# m1_32818_24542# vss nfet$221
Xnfet$214_6 m1_n1133_19550# m1_n1133_19550# vss vss m1_n695_20470# vss nfet$214
Xnfet$216_16 m1_26873_21786# vss m1_27003_21590# vss nfet$216
Xnfet$232_15 m1_17697_15478# m1_17697_15478# m1_n2543_20130# m1_n2543_20130# m1_20407_20470#
+ vss nfet$232
Xpfet$204_11 vdd vdd m1_32817_25662# m1_32675_25947# pfet$204
Xnfet$212_3 m1_488_21786# vss m1_2912_25858# vss nfet$212
Xpfet$204_4 vdd vdd m1_488_21786# m1_n789_25858# pfet$204
Xnfet$213_17 m1_12935_21590# m1_12935_21590# m1_14422_22513# m1_14422_22513# m1_13394_21586#
+ vss nfet$213
Xpfet$196_91 vdd vdd m1_23356_21786# pd8 pfet$196
Xpfet$196_80 vdd vdd m1_17058_24346# m1_n7513_20152# pfet$196
Xpfet$202_1 vdd vdd m1_4620_20152# m1_n3218_15478# pfet$202
Xpfet$201_12 vdd vdd m1_26676_16080# m1_n7513_20152# pfet$201
Xnfet$239_8 m1_n4623_25487# vss m1_n4464_25980# vss nfet$239
Xnfet$224_16 m1_28624_21786# m1_28624_21786# vss vss m1_27462_21586# vss nfet$224
Xpfet$198_26 vdd vdd vdd m1_16911_22102# m1_16452_21590# m1_16452_21590# pfet$198
Xpfet$198_15 vdd m1_354_22513# m1_354_22513# m1_n46_22402# m1_488_21786# m1_488_21786#
+ pfet$198
Xnfet$228_1 m1_30256_19792# vss m1_32818_20470# vss nfet$228
Xnfet$235_2 m1_n6788_16080# m1_n6788_16080# m1_n7247_17714# m1_n7247_17714# m1_n6690_16398#
+ vss nfet$235
Xnfet$214_7 m1_n7383_17599# m1_n7383_17599# vss vss m1_n63_20470# vss nfet$214
Xnfet$216_17 m1_25107_21786# vss m1_25739_21786# vss nfet$216
Xnfet$232_16 m1_25722_20152# m1_25722_20152# m1_n3206_20274# m1_n3206_20274# m1_24556_20470#
+ vss nfet$232
Xpfet$225_0 vdd m1_n6380_21786# m1_n6380_21786# m1_n5019_19550# m1_n5227_20152# m1_n5227_20152#
+ pfet$225
Xnfet$240_0 m1_n9952_24224# m1_n9952_24224# m1_n10308_24542# m1_n10308_24542# m1_n9854_24542#
+ vss nfet$240
Xpfet$204_12 vdd vdd m1_32193_25858# m1_25107_21786# pfet$204
Xpfet$204_5 vdd vdd m1_326_24346# m1_n7513_20152# pfet$204
Xnfet$212_4 m1_2912_25858# vss m1_3049_25662# vss nfet$212
Xpfet$196_92 vdd vdd m1_28492_25858# m1_29607_24346# pfet$196
Xpfet$196_81 vdd vdd m1_18339_24542# m1_15943_25858# pfet$196
Xpfet$196_70 vdd vdd m1_14156_24542# m1_11760_25858# pfet$196
Xpfet$202_2 vdd vdd m1_1103_20152# m1_n7401_15478# pfet$202
Xpfet$201_13 vdd vdd m1_25747_17714# m1_26217_17714# pfet$201
Xnfet$239_9 m1_n3184_24224# vss m1_n3541_23922# vss nfet$239
Xnfet$224_17 m1_29256_21786# m1_29256_21786# vss vss m1_28094_21586# vss nfet$224
Xpfet$198_27 vdd m1_14422_22513# m1_14422_22513# m1_14022_22402# m1_14556_21786# m1_14556_21786#
+ pfet$198
Xpfet$198_16 vdd m1_24973_22513# m1_24973_22513# m1_23945_22102# m1_25739_21786# m1_25739_21786#
+ pfet$198
Xnfet$228_2 m1_31535_19792# m1_32818_20470# vss vss nfet$228
Xnfet$235_3 m1_n6172_16202# m1_n6172_16202# vss vss m1_n6690_16398# vss nfet$235
Xnfet$214_8 m1_27003_19550# m1_27003_19550# vss vss m1_27441_20470# vss nfet$214
Xnfet$232_17 m1_21880_15478# m1_21880_15478# m1_n3206_20274# m1_n3206_20274# m1_23924_20470#
+ vss nfet$232
Xnfet$233_0 m1_35837_22102# vss m1_n7513_20152# vss nfet$233
Xnfet$240_1 m1_n9336_24346# m1_n9336_24346# m1_n8625_26174# m1_n8625_26174# m1_n8389_25502#
+ vss nfet$240
Xpfet$225_1 vdd vdd vdd m1_n5019_22344# m1_n4485_21904# m1_n4485_21904# pfet$225
Xpfet$218_0 vdd m1_n10309_25662# m1_n10572_23922# m1_n10796_25662# pfet$218
Xpfet$204_13 vdd vdd m1_33790_24346# m1_n7513_20152# pfet$204
Xnfet$212_5 m1_2912_25858# m1_3536_25662# m1_3273_23922# vss nfet$212
Xpfet$204_6 vdd vdd m1_n290_24224# m1_n910_23922# pfet$204
Xpfet$196_93 vdd m1_28991_24224# m1_30095_25658# m1_28010_25858# pfet$196
Xpfet$196_82 vdd vdd m1_21241_24346# m1_n7513_20152# pfet$196
Xpfet$196_71 vdd vdd m1_11039_21786# m1_11760_25858# pfet$196
Xpfet$196_60 vdd vdd m1_20126_25858# m1_21241_24346# pfet$196
Xpfet$202_3 vdd vdd m1_5901_19550# m1_649_17714# pfet$202
Xpfet$200_0 vdd vdd m1_n1133_21590# m1_n1263_21786# pfet$200
Xpfet$198_28 vdd m1_14422_22513# m1_14422_22513# m1_13394_22102# m1_15188_21786# m1_15188_21786#
+ pfet$198
Xpfet$198_17 vdd m1_21456_22513# m1_21456_22513# m1_21056_22402# m1_21590_21786# m1_21590_21786#
+ pfet$198
Xnfet$235_4 m1_28113_15778# m1_28113_15778# m1_28003_18030# m1_28003_18030# m1_28239_17358#
+ vss nfet$235
Xnfet$228_3 m1_30256_22102# vss m1_32818_21586# vss nfet$228
Xnfet$214_9 m1_25747_17714# m1_25747_17714# vss vss m1_28073_20470# vss nfet$214
Xpfet$198_0 vdd vdd vdd m1_n674_22102# m1_n1133_21590# m1_n1133_21590# pfet$198
Xnfet$226_0 m1_34843_21786# m1_34843_21786# m1_34093_22102# m1_34093_22102# m1_34329_21430#
+ vss nfet$226
Xnfet$240_2 m1_n8848_25658# m1_n8848_25658# vss vss m1_n8389_25502# vss nfet$240
Xpfet$225_2 vdd m1_n5764_21786# m1_n5764_21786# m1_n5019_22344# m1_n5227_21418# m1_n5227_21418#
+ pfet$225
Xpfet$218_1 vdd m1_n9952_24224# m1_n8848_25658# m1_n10933_25858# pfet$218
Xnfet$212_6 m1_3049_25662# m1_3893_24224# m1_4997_25658# vss nfet$212
Xpfet$204_7 vdd vdd m1_32330_25662# m1_32193_25858# pfet$204
Xpfet$196_94 vdd m1_28492_25858# vdd m1_30095_25658# pfet$196
Xpfet$196_83 vdd m1_21729_25658# m1_22522_24542# m1_19781_25662# pfet$196
Xpfet$196_72 vdd m1_13363_25658# m1_14156_24542# m1_11415_25662# pfet$196
Xpfet$196_61 vdd m1_24452_24542# vdd m1_25424_24346# pfet$196
Xpfet$196_50 vdd vdd m1_20268_25662# m1_20126_25858# pfet$196
Xpfet$202_4 vdd vdd m1_12935_19550# m1_9015_17714# pfet$202
Xpfet$200_1 vdd vdd m1_11671_21786# m1_11039_21786# pfet$200
Xpfet$198_29 vdd vdd vdd m1_14022_22402# m1_12805_21786# m1_12805_21786# pfet$198
Xpfet$198_18 vdd vdd vdd m1_24573_22402# m1_23356_21786# m1_23356_21786# pfet$198
Xnfet$235_5 m1_26676_16080# m1_26676_16080# vss vss m1_28239_17358# vss nfet$235
Xnfet$211_20 m1_21241_24346# m1_21241_24346# m1_20126_25858# m1_20126_25858# m1_22188_25502#
+ vss nfet$211
Xpfet$198_1 vdd m1_7388_22513# m1_7388_22513# m1_6988_22402# m1_7522_21786# m1_7522_21786#
+ pfet$198
Xnfet$226_1 m1_28490_22513# m1_28490_22513# vss vss m1_34329_21430# vss nfet$226
Xnfet$219_0 m1_n3534_17714# vss m1_n6433_17343# vss nfet$219
Xnfet$240_3 m1_n9336_24346# m1_n9336_24346# vss vss m1_n9854_24542# vss nfet$240
Xpfet$218_2 vdd m1_n4362_24346# m1_n4847_25662# m1_n4464_25980# pfet$218
Xnfet$212_7 m1_3049_25662# m1_3273_23922# m1_3537_24542# vss nfet$212
Xpfet$204_8 vdd vdd m1_33174_24224# m1_32554_23922# pfet$204
Xpfet$196_95 vdd vdd m1_28991_24224# m1_28371_23922# pfet$196
Xpfet$196_84 vdd vdd m1_23827_25858# m1_18073_21786# pfet$196
Xpfet$196_73 vdd m1_16086_24542# vdd m1_17058_24346# pfet$196
Xpfet$196_62 vdd vdd m1_24452_24542# m1_24808_24224# pfet$196
Xpfet$196_51 vdd vdd m1_20625_24224# m1_20005_23922# pfet$196
Xpfet$196_40 vdd vdd m1_11760_25858# m1_12875_24346# pfet$196
Xpfet$223_0 vdd vdd m1_n7186_25858# m1_n10452_25858# pfet$223
Xpfet$202_5 vdd vdd m1_8137_20152# m1_965_15478# pfet$202
Xpfet$200_2 vdd vdd m1_12935_21590# m1_12805_21786# pfet$200
Xpfet$198_19 vdd m1_24973_22513# m1_24973_22513# m1_24573_22402# m1_25107_21786# m1_25107_21786#
+ pfet$198
Xnfet$235_6 m1_27292_16202# m1_27292_16202# vss vss m1_26774_16398# vss nfet$235
Xnfet$211_21 m1_28991_24224# m1_28991_24224# m1_28635_24542# m1_28635_24542# m1_29089_24542#
+ vss nfet$211
Xnfet$211_10 m1_17546_25658# m1_17546_25658# vss vss m1_18005_25502# vss nfet$211
Xpfet$198_2 vdd m1_7388_22513# m1_7388_22513# m1_6360_22102# m1_8154_21786# m1_8154_21786#
+ pfet$198
Xnfet$240_4 m1_n4978_24224# m1_n4978_24224# m1_n10452_25858# m1_n10452_25858# m1_n4880_24542#
+ vss nfet$240
Xnfet$226_2 m1_9645_21447# m1_9645_21447# vss vss m1_30492_21430# vss nfet$226
Xnfet$219_1 m1_n7513_20152# vss m1_n6788_16080# vss nfet$219
Xpfet$218_3 vdd m1_n3184_24224# m1_n3651_26174# m1_n4623_25487# pfet$218
Xnfet$212_8 m1_3394_25858# vss m1_3536_25662# vss nfet$212
Xpfet$204_9 vdd vdd m1_28624_21786# m1_32675_25947# pfet$204
Xnfet$231_0 m1_7198_15778# m1_7198_15778# m1_7088_18030# m1_7088_18030# m1_7324_17358#
+ vss nfet$231
Xpfet$196_41 vdd vdd m1_9288_21786# pd4 pfet$196
Xpfet$216_0 vdd vdd m1_n7513_20152# m1_35837_22102# pfet$216
Xpfet$196_30 vdd vdd m1_2912_25858# m1_488_21786# pfet$196
Xpfet$223_1 vdd m1_n7186_25858# vdd m1_n6111_25858# pfet$223
Xpfet$196_96 vdd m1_28635_24542# vdd m1_29607_24346# pfet$196
Xpfet$196_85 vdd m1_24188_23922# m1_24452_24542# m1_23827_25858# pfet$196
Xpfet$196_74 vdd vdd m1_14556_21786# m1_15943_25858# pfet$196
Xpfet$196_63 vdd vdd m1_19781_25662# m1_19644_25858# pfet$196
Xpfet$196_52 vdd m1_20268_25662# m1_20005_23922# m1_19781_25662# pfet$196
Xpfet$202_6 vdd vdd m1_9418_19550# m1_4832_17714# pfet$202
Xpfet$200_3 vdd vdd m1_9418_21590# m1_9288_21786# pfet$200
Xnfet$214_10 m1_9015_17714# m1_9015_17714# vss vss m1_14005_20470# vss nfet$214
Xnfet$235_7 m1_26676_16080# m1_26676_16080# m1_26217_17714# m1_26217_17714# m1_26774_16398#
+ vss nfet$235
Xnfet$211_22 m1_29607_24346# m1_29607_24346# vss vss m1_29089_24542# vss nfet$211
Xnfet$211_11 m1_16442_24224# m1_16442_24224# m1_16086_24542# m1_16086_24542# m1_16540_24542#
+ vss nfet$211
Xpfet$198_3 vdd m1_9645_21447# m1_9645_21447# m1_10505_22402# m1_11039_21786# m1_11039_21786#
+ pfet$198
Xpfet$199_30 vdd vdd vdd m1_24560_19550# m1_21880_15478# m1_21880_15478# pfet$199
Xnfet$226_3 m1_7388_22513# m1_7388_22513# m1_30256_22102# m1_30256_22102# m1_30492_21430#
+ vss nfet$226
Xnfet$219_2 m1_n4994_16080# vss m1_n5351_15778# vss nfet$219
Xnfet$240_5 m1_n4362_24346# m1_n4362_24346# vss vss m1_n4880_24542# vss nfet$240
Xpfet$218_4 vdd m1_n2567_23922# m1_n3184_24224# m1_n4464_25980# pfet$218
Xpfet$196_0 vdd vdd m1_3049_25662# m1_2912_25858# pfet$196
Xnfet$212_9 m1_3273_23922# vss m1_3893_24224# vss nfet$212
Xnfet$231_1 m1_5761_16080# m1_5761_16080# vss vss m1_7324_17358# vss nfet$231
Xnfet$224_0 m1_11039_21786# m1_11039_21786# vss vss m1_9877_21586# vss nfet$224
Xnfet$217_10 m1_26063_15478# vss m1_29239_20152# vss nfet$217
Xpfet$209_0 vdd vdd m1_n1263_21786# pd1 pfet$209
Xpfet$196_97 vdd vdd m1_21590_21786# m1_24309_25858# pfet$196
Xpfet$196_86 vdd m1_28634_25662# m1_28371_23922# m1_28147_25662# pfet$196
Xpfet$196_75 vdd vdd m1_19644_25858# m1_14556_21786# pfet$196
Xpfet$196_64 vdd vdd m1_22522_24542# m1_20126_25858# pfet$196
Xpfet$196_53 vdd m1_20625_24224# m1_21729_25658# m1_19644_25858# pfet$196
Xpfet$196_42 vdd m1_11760_25858# vdd m1_13363_25658# pfet$196
Xpfet$196_31 vdd m1_3273_23922# m1_3537_24542# m1_2912_25858# pfet$196
Xpfet$196_20 vdd vdd m1_4509_24346# m1_n7513_20152# pfet$196
Xpfet$202_7 vdd vdd m1_11654_20152# m1_5148_15478# pfet$202
Xnfet$214_11 m1_13198_17714# m1_13198_17714# vss vss m1_17522_20470# vss nfet$214
Xpfet$200_4 vdd vdd m1_8154_21786# m1_7522_21786# pfet$200
Xpfet$198_4 vdd vdd vdd m1_9877_22102# m1_9418_21590# m1_9418_21590# pfet$198
Xnfet$211_23 m1_25424_24346# m1_25424_24346# m1_24309_25858# m1_24309_25858# m1_26371_25502#
+ vss nfet$211
Xnfet$211_12 m1_17058_24346# m1_17058_24346# m1_15943_25858# m1_15943_25858# m1_18005_25502#
+ vss nfet$211
Xpfet$199_31 vdd m1_n2543_20130# m1_n2543_20130# m1_20407_19850# m1_19969_19550# m1_19969_19550#
+ pfet$199
Xpfet$199_20 vdd m1_n3822_21786# m1_n3822_21786# m1_14009_19550# m1_9015_17714# m1_9015_17714#
+ pfet$199
Xnfet$219_3 m1_n6433_17343# vss m1_n6274_17836# vss nfet$219
Xnfet$240_6 m1_n4978_24224# m1_n4978_24224# vss vss m1_n3415_25502# vss nfet$240
Xpfet$196_1 vdd m1_3536_25662# m1_3273_23922# m1_3049_25662# pfet$196
Xpfet$218_5 vdd m1_n10572_23922# m1_n10308_24542# m1_n10933_25858# pfet$218
Xpfet$209_1 vdd vdd m1_2254_21786# pd2 pfet$209
Xnfet$217_0 m1_n3534_17714# vss m1_2384_19550# vss nfet$217
Xnfet$231_2 m1_9944_16080# m1_9944_16080# vss vss m1_11507_17358# vss nfet$231
Xnfet$224_1 m1_11671_21786# m1_11671_21786# vss vss m1_10509_21586# vss nfet$224
Xpfet$196_98 vdd m1_30095_25658# m1_30888_24542# m1_28147_25662# pfet$196
Xpfet$196_87 vdd vdd m1_28147_25662# m1_28010_25858# pfet$196
Xpfet$196_76 vdd m1_20005_23922# m1_20269_24542# m1_19644_25858# pfet$196
Xpfet$196_65 vdd vdd m1_18073_21786# m1_20126_25858# pfet$196
Xpfet$196_54 vdd vdd m1_24808_24224# m1_24188_23922# pfet$196
Xpfet$196_43 vdd vdd m1_12805_21786# pd5 pfet$196
Xnfet$217_11 m1_9331_15478# vss m1_15171_20152# vss nfet$217
Xpfet$196_32 vdd vdd m1_7720_24542# m1_8076_24224# pfet$196
Xpfet$196_21 vdd m1_7456_23922# m1_7720_24542# m1_7095_25858# pfet$196
Xpfet$196_10 vdd m1_8076_24224# m1_9180_25658# m1_7095_25858# pfet$196
Xpfet$202_8 vdd vdd m1_n1133_19550# m1_n7383_17599# pfet$202
Xpfet$221_0 vdd vdd m1_n4485_20152# m1_n3822_20130# pfet$221
Xnfet$214_12 m1_16452_19550# m1_16452_19550# vss vss m1_16890_20470# vss nfet$214
Xpfet$200_5 vdd vdd m1_1120_21786# m1_488_21786# pfet$200
Xnfet$247_0 m1_n6839_20152# vss m1_n8145_21908# vss nfet$247
Xnfet$211_24 m1_30095_25658# m1_30095_25658# vss vss m1_30554_25502# vss nfet$211
Xnfet$211_13 m1_13363_25658# m1_13363_25658# vss vss m1_13822_25502# vss nfet$211
Xpfet$199_32 vdd m1_n2543_20130# m1_n2543_20130# m1_21043_19550# m1_17381_17714# m1_17381_17714#
+ pfet$199
Xpfet$199_21 vdd vdd vdd m1_13373_19850# m1_15171_20152# m1_15171_20152# pfet$199
Xpfet$199_10 vdd vdd vdd m1_9856_19850# m1_11654_20152# m1_11654_20152# pfet$199
Xpfet$198_5 vdd m1_9645_21447# m1_9645_21447# m1_9877_22102# m1_11671_21786# m1_11671_21786#
+ pfet$198
Xnfet$219_4 m1_n7247_17714# vss m1_n4377_15778# vss nfet$219
Xnfet$240_7 m1_n3541_23922# m1_n3541_23922# m1_n3651_26174# m1_n3651_26174# m1_n3415_25502#
+ vss nfet$240
Xpfet$196_2 vdd vdd m1_3394_25858# m1_4509_24346# pfet$196
Xpfet$218_6 vdd m1_n8848_25658# m1_n8055_24542# m1_n10796_25662# pfet$218
Xnfet$217_1 m1_n3218_15478# vss m1_4620_20152# vss nfet$217
Xnfet$231_3 m1_11381_15778# m1_11381_15778# m1_11271_18030# m1_11271_18030# m1_11507_17358#
+ vss nfet$231
Xnfet$224_2 m1_8154_21786# m1_8154_21786# vss vss m1_6992_21586# vss nfet$224
Xpfet$196_99 vdd vdd m1_26705_24542# m1_24309_25858# pfet$196
Xpfet$209_2 vdd vdd m1_26873_21786# pd9 pfet$209
Xpfet$196_88 vdd vdd m1_28634_25662# m1_28492_25858# pfet$196
Xpfet$196_77 vdd vdd m1_20269_24542# m1_20625_24224# pfet$196
Xpfet$196_66 vdd vdd m1_15461_25858# m1_11039_21786# pfet$196
Xpfet$196_55 vdd m1_24451_25662# m1_24188_23922# m1_23964_25662# pfet$196
Xpfet$196_44 vdd m1_15943_25858# vdd m1_17546_25658# pfet$196
Xnfet$217_12 m1_13514_15478# vss m1_18688_20152# vss nfet$217
Xpfet$196_33 vdd vdd m1_7522_21786# m1_7577_25858# pfet$196
Xpfet$196_22 vdd vdd m1_3537_24542# m1_3893_24224# pfet$196
Xpfet$196_11 vdd vdd m1_7719_25662# m1_7577_25858# pfet$196
Xpfet$202_9 vdd vdd m1_27003_19550# m1_25747_17714# pfet$202
Xpfet$214_0 vdd vdd m1_n7247_17714# m1_n6788_16080# pfet$214
Xpfet$221_1 vdd m1_n4485_21904# vdd m1_9624_19404# pfet$221
Xnfet$214_13 m1_19969_19550# m1_19969_19550# vss vss m1_20407_20470# vss nfet$214
Xpfet$200_6 vdd vdd m1_5901_21590# m1_5771_21786# pfet$200
Xnfet$239_10 vss vss m1_n4978_24224# vss nfet$239
Xnfet$211_25 m1_29607_24346# m1_29607_24346# m1_28492_25858# m1_28492_25858# m1_30554_25502#
+ vss nfet$211
Xnfet$211_14 m1_12875_24346# m1_12875_24346# m1_11760_25858# m1_11760_25858# m1_13822_25502#
+ vss nfet$211
Xpfet$198_6 vdd vdd vdd m1_10505_22402# m1_9288_21786# m1_9288_21786# pfet$198
Xpfet$199_33 vdd m1_n3206_20274# m1_n3206_20274# m1_24560_19550# m1_21564_17714# m1_21564_17714#
+ pfet$199
Xpfet$199_22 vdd vdd vdd m1_14009_19550# m1_9331_15478# m1_9331_15478# pfet$199
Xpfet$199_11 vdd vdd vdd m1_10492_19550# m1_5148_15478# m1_5148_15478# pfet$199
Xnfet$219_5 m1_n7247_17714# vss m1_n6657_17518# vss nfet$219
Xpfet$196_3 vdd m1_3394_25858# vdd m1_4997_25658# pfet$196
Xpfet$218_7 vdd m1_n3541_23922# m1_n4362_24346# m1_n4623_25487# pfet$218
Xnfet$217_2 m1_n7401_15478# vss m1_1103_20152# vss nfet$217
Xnfet$231_4 m1_10560_16202# m1_10560_16202# vss vss m1_10042_16398# vss nfet$231
Xnfet$224_3 m1_7522_21786# m1_7522_21786# vss vss m1_6360_21586# vss nfet$224
Xpfet$196_89 vdd vdd m1_19839_21786# pd7 pfet$196
Xpfet$196_78 vdd m1_20269_24542# vdd m1_21241_24346# pfet$196
Xpfet$196_67 vdd m1_15822_23922# m1_16086_24542# m1_15461_25858# pfet$196
Xpfet$196_56 vdd m1_24808_24224# m1_25912_25658# m1_23827_25858# pfet$196
Xpfet$196_45 vdd vdd m1_16442_24224# m1_15822_23922# pfet$196
Xnfet$217_13 m1_13198_17714# vss m1_16452_19550# vss nfet$217
Xpfet$196_34 vdd m1_9180_25658# m1_9973_24542# m1_7232_25662# pfet$196
Xpfet$196_23 vdd m1_3537_24542# vdd m1_4509_24346# pfet$196
Xpfet$196_12 vdd m1_7577_25858# vdd m1_9180_25658# pfet$196
Xpfet$207_0 vdd m1_31535_19792# vdd m1_17939_22513# pfet$207
Xnfet$222_0 pd1 vss m1_n1263_21786# vss nfet$222
Xpfet$214_1 vdd m1_n7247_17714# vdd m1_n6172_16202# pfet$214
Xpfet$221_2 vdd m1_n5227_21418# vdd m1_2590_19404# pfet$221
Xpfet$200_7 vdd vdd m1_4637_21786# m1_4005_21786# pfet$200
Xnfet$214_14 m1_17381_17714# m1_17381_17714# vss vss m1_21039_20470# vss nfet$214
Xnfet$239_11 m1_n10452_25858# vss m1_n4847_25662# vss nfet$239
Xpfet$197_110 vdd vdd m1_10458_17836# m1_10299_17343# pfet$197
Xnfet$211_26 m1_25912_25658# m1_25912_25658# vss vss m1_26371_25502# vss nfet$211
Xnfet$211_15 m1_25424_24346# m1_25424_24346# vss vss m1_24906_24542# vss nfet$211
Xpfet$198_7 vdd m1_354_22513# m1_354_22513# m1_n674_22102# m1_1120_21786# m1_1120_21786#
+ pfet$198
Xpfet$199_34 vdd m1_n3206_20274# m1_n3206_20274# m1_23924_19850# m1_23486_19550# m1_23486_19550#
+ pfet$199
Xpfet$199_23 vdd vdd vdd m1_16890_19850# m1_18688_20152# m1_18688_20152# pfet$199
Xpfet$199_12 vdd m1_6107_19404# m1_6107_19404# m1_6975_19550# m1_649_17714# m1_649_17714#
+ pfet$199
Xnfet$219_6 m1_n7247_17714# vss m1_n7383_17599# vss nfet$219
Xpfet$196_4 vdd vdd m1_3893_24224# m1_3273_23922# pfet$196
Xnfet$212_80 m1_28147_25662# m1_28991_24224# m1_30095_25658# vss nfet$212
Xnfet$217_3 m1_649_17714# vss m1_5901_19550# vss nfet$217
Xnfet$231_5 m1_9944_16080# m1_9944_16080# m1_9485_17714# m1_9485_17714# m1_10042_16398#
+ vss nfet$231
Xnfet$224_4 m1_1120_21786# m1_1120_21786# vss vss m1_n42_21586# vss nfet$224
Xpfet$196_57 vdd vdd m1_24451_25662# m1_24309_25858# pfet$196
Xpfet$196_46 vdd m1_16442_24224# m1_17546_25658# m1_15461_25858# pfet$196
Xnfet$217_14 m1_21564_17714# vss m1_23486_19550# vss nfet$217
Xpfet$196_35 vdd m1_7720_24542# vdd m1_8692_24346# pfet$196
Xpfet$196_24 vdd vdd m1_5790_24542# m1_3394_25858# pfet$196
Xpfet$196_13 vdd vdd m1_12259_24224# m1_11639_23922# pfet$196
Xpfet$196_79 vdd m1_17546_25658# m1_18339_24542# m1_15598_25662# pfet$196
Xpfet$196_68 vdd vdd m1_16086_24542# m1_16442_24224# pfet$196
Xnfet$222_1 pd2 vss m1_2254_21786# vss nfet$222
Xnfet$215_0 m1_9485_17714# vss m1_9015_17714# vss nfet$215
Xpfet$207_1 vdd vdd m1_30256_19792# m1_21456_22513# pfet$207
Xpfet$214_2 vdd vdd m1_n5461_18030# m1_n5351_15778# pfet$214
Xpfet$221_3 vdd vdd m1_n5227_21418# m1_6107_19404# pfet$221
Xpfet$200_8 vdd vdd m1_2384_21590# m1_2254_21786# pfet$200
Xnfet$214_15 m1_21564_17714# m1_21564_17714# vss vss m1_24556_20470# vss nfet$214
Xnfet$239_12 m1_n10452_25858# vss m1_n5571_25662# vss nfet$239
Xpfet$202_10 vdd vdd m1_29239_20152# m1_26063_15478# pfet$202
Xpfet$197_100 vdd vdd m1_23820_18030# m1_23930_15778# pfet$197
Xnfet$215_80 m1_18824_17836# m1_19747_15778# m1_18926_16202# vss nfet$215
Xnfet$211_27 m1_12875_24346# m1_12875_24346# vss vss m1_12357_24542# vss nfet$211
Xnfet$211_16 m1_24808_24224# m1_24808_24224# m1_24452_24542# m1_24452_24542# m1_24906_24542#
+ vss nfet$211
Xpfet$198_8 vdd vdd vdd m1_6360_22102# m1_5901_21590# m1_5901_21590# pfet$198
Xpfet$199_35 vdd m1_n3822_21786# m1_n3822_21786# m1_13373_19850# m1_12935_19550# m1_12935_19550#
+ pfet$199
Xpfet$199_24 vdd m1_n1927_20274# m1_n1927_20274# m1_16890_19850# m1_16452_19550# m1_16452_19550#
+ pfet$199
Xpfet$199_13 vdd m1_n927_19404# m1_n927_19404# m1_n695_19850# m1_n1133_19550# m1_n1133_19550#
+ pfet$199
Xnfet$219_7 m1_26217_17714# vss m1_26807_17518# vss nfet$219
Xnfet$245_0 m1_n927_19404# m1_n927_19404# vss vss m1_n6282_20470# vss nfet$245
Xpfet$196_5 vdd m1_3893_24224# m1_4997_25658# m1_2912_25858# pfet$196
Xnfet$212_81 m1_n7513_20152# vss m1_25424_24346# vss nfet$212
Xnfet$212_70 m1_21590_21786# vss m1_28010_25858# vss nfet$212
Xnfet$217_4 m1_4832_17714# vss m1_9418_19550# vss nfet$217
Xnfet$231_6 m1_1578_16080# m1_1578_16080# vss vss m1_3141_17358# vss nfet$231
Xnfet$224_5 m1_4005_21786# m1_4005_21786# vss vss m1_2843_21586# vss nfet$224
Xnfet$217_15 m1_17697_15478# vss m1_22205_20152# vss nfet$217
Xpfet$196_69 vdd vdd m1_12875_24346# m1_n7513_20152# pfet$196
Xpfet$196_58 vdd vdd m1_23964_25662# m1_23827_25858# pfet$196
Xpfet$196_47 vdd vdd m1_15943_25858# m1_17058_24346# pfet$196
Xpfet$196_36 vdd vdd m1_8692_24346# m1_n7513_20152# pfet$196
Xpfet$196_25 vdd vdd m1_4005_21786# m1_3394_25858# pfet$196
Xpfet$196_14 vdd vdd m1_11902_25662# m1_11760_25858# pfet$196
Xnfet$222_2 pd9 vss m1_26873_21786# vss nfet$222
Xnfet$215_1 m1_9015_17714# vss m1_6116_17343# vss nfet$215
Xpfet$207_2 vdd m1_30256_19792# vdd m1_24973_22513# pfet$207
Xpfet$214_3 vdd m1_n5461_18030# vdd m1_n6788_16080# pfet$214
Xpfet$221_4 vdd vdd m1_n4485_21904# m1_n3822_21786# pfet$221
Xpfet$197_90 vdd m1_19747_15778# m1_18926_16202# m1_18665_17343# pfet$197
Xpfet$212_0 vdd vdd fout m1_34093_22102# pfet$212
Xpfet$200_9 vdd vdd m1_22222_21786# m1_21590_21786# pfet$200
Xnfet$214_16 m1_23486_19550# m1_23486_19550# vss vss m1_23924_20470# vss nfet$214
Xnfet$239_13 fin vss m1_n4623_25487# vss nfet$239
Xpfet$197_101 vdd vdd m1_19637_18030# m1_19747_15778# pfet$197
Xpfet$202_11 vdd vdd m1_18688_20152# m1_13514_15478# pfet$202
Xnfet$215_81 m1_13198_17714# vss m1_10299_17343# vss nfet$215
Xnfet$215_70 m1_n7513_20152# vss m1_18310_16080# vss nfet$215
Xpfet$198_9 vdd m1_3871_22513# m1_3871_22513# m1_3471_22402# m1_4005_21786# m1_4005_21786#
+ pfet$198
Xnfet$211_17 m1_20625_24224# m1_20625_24224# m1_20269_24542# m1_20269_24542# m1_20723_24542#
+ vss nfet$211
Xpfet$199_25 vdd vdd vdd m1_17526_19550# m1_13514_15478# m1_13514_15478# pfet$199
Xpfet$199_14 vdd m1_n927_19404# m1_n927_19404# m1_n59_19550# m1_n7383_17599# m1_n7383_17599#
+ pfet$199
Xnfet$219_8 m1_n7513_20152# vss m1_26676_16080# vss nfet$219
Xpfet$196_6 vdd vdd m1_3536_25662# m1_3394_25858# pfet$196
Xnfet$238_0 m1_n3822_20130# m1_n3822_20130# m1_n4485_20152# m1_n4485_20152# m1_n3724_20470#
+ vss nfet$238
Xnfet$245_1 m1_n2543_20130# m1_n2543_20130# m1_n5227_20152# m1_n5227_20152# m1_n2445_20470#
+ vss nfet$245
Xnfet$212_82 m1_11415_25662# m1_12259_24224# m1_13363_25658# vss nfet$212
Xnfet$212_71 m1_28147_25662# m1_28371_23922# m1_28635_24542# vss nfet$212
Xnfet$212_60 pd6 vss m1_16322_21786# vss nfet$212
Xnfet$217_5 m1_965_15478# vss m1_8137_20152# vss nfet$217
Xnfet$231_7 m1_5761_16080# m1_5761_16080# m1_5302_17714# m1_5302_17714# m1_5859_16398#
+ vss nfet$231
Xnfet$224_6 m1_4637_21786# m1_4637_21786# vss vss m1_3475_21586# vss nfet$224
Xpfet$196_59 vdd vdd m1_16322_21786# pd6 pfet$196
Xpfet$196_48 vdd m1_16085_25662# m1_15822_23922# m1_15598_25662# pfet$196
Xnfet$217_16 m1_17381_17714# vss m1_19969_19550# vss nfet$217
Xpfet$196_37 vdd vdd m1_9973_24542# m1_7577_25858# pfet$196
Xpfet$196_26 vdd m1_4997_25658# m1_5790_24542# m1_3049_25662# pfet$196
Xpfet$196_15 vdd m1_11902_25662# m1_11639_23922# m1_11415_25662# pfet$196
Xnfet$215_2 m1_6275_17836# m1_7555_16080# m1_7088_18030# vss nfet$215
Xpfet$207_3 vdd vdd m1_34843_21786# m1_34093_19792# pfet$207
Xpfet$214_4 vdd vdd m1_26217_17714# m1_26676_16080# pfet$214
Xpfet$221_5 vdd m1_n6839_21786# vdd m1_n5764_21786# pfet$221
Xpfet$197_91 vdd m1_24287_16080# m1_23820_18030# m1_22848_17343# pfet$197
Xpfet$197_80 vdd vdd m1_15564_15778# m1_15921_16080# pfet$197
Xnfet$214_17 m1_12935_19550# m1_12935_19550# vss vss m1_13373_20470# vss nfet$214
Xnfet$220_0 m1_n10452_25858# vss m1_n1271_25858# vss nfet$220
Xpfet$205_0 vdd vdd m1_n646_24542# m1_n290_24224# pfet$205
Xpfet$202_12 vdd vdd m1_15171_20152# m1_9331_15478# pfet$202
Xpfet$197_102 vdd vdd m1_13198_17714# m1_13668_17714# pfet$197
Xnfet$215_82 m1_10299_17343# vss m1_10458_17836# vss nfet$215
Xnfet$215_71 m1_14641_17836# m1_15921_16080# m1_15454_18030# vss nfet$215
Xnfet$215_60 m1_18665_17343# vss m1_18824_17836# vss nfet$215
Xnfet$211_18 m1_21241_24346# m1_21241_24346# vss vss m1_20723_24542# vss nfet$211
Xpfet$199_26 vdd m1_n1927_20274# m1_n1927_20274# m1_17526_19550# m1_13198_17714# m1_13198_17714#
+ pfet$199
Xpfet$199_15 vdd vdd vdd m1_n59_19550# m1_n7401_15478# m1_n7401_15478# pfet$199
Xnfet$219_9 m1_n10452_25858# vss m1_27031_17343# vss nfet$219
.ends

.subckt asc_drive_buffer$4 vss in vdd out
Xpfet$265_0 vdd vdd m1_3466_n454# in pfet$265
Xpfet$263_0 m1_4274_n1060# vdd vdd m1_4274_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ vdd m1_4002_n1060# m1_4002_n1060# pfet$263
Xnfet$283_0 m1_3466_n454# vss m1_4002_n1060# vss nfet$283
Xnfet$281_0 m1_4274_n1060# vss m1_4002_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ m1_4274_n1060# vss m1_4002_n1060# vss nfet$281
Xpfet$264_0 vdd vdd m1_4002_n1060# m1_3466_n454# pfet$264
Xpfet$262_0 out out m1_4274_n1060# vdd m1_4274_n1060# out vdd vdd m1_4274_n1060# out
+ m1_4274_n1060# m1_4274_n1060# out m1_4274_n1060# vdd m1_4274_n1060# vdd m1_4274_n1060#
+ pfet$262
Xnfet$284_0 in vss m1_3466_n454# vss nfet$284
Xnfet$282_0 out out vss m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# m1_4274_n1060#
+ m1_4274_n1060# out m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# vss vss
+ nfet$282
.ends

.subckt pfet$275 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$298 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$267 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$272 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$270 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$296 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt nfet$289 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$294 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$287 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$277 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt nfet$292 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$285 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$290 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt pfet$268 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$273 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$266 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$271 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt nfet$297 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt nfet$295 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$288 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$278 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$293 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt nfet$286 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$291 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$276 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt pfet$269 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$274 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt asc_PFD_DFF_20250831 vss fref down up vdd fdiv
Xpfet$275_17 vdd vdd m1_n5649_n11124# m1_n5867_n10544# pfet$275
Xnfet$298_0 up up m1_5895_n8089# m1_5895_n8089# m1_5043_n9245# vss nfet$298
Xpfet$267_3 vdd vdd m1_2779_n3533# m1_2068_n5361# pfet$267
Xpfet$275_18 vdd vdd m1_n5867_n10544# fdiv pfet$275
Xpfet$272_1 vdd vdd m1_n5650_n4045# m1_n5868_n3849# pfet$272
Xnfet$298_1 down down vss vss m1_5043_n9245# vss nfet$298
Xpfet$272_2 vdd vdd m1_n3885_n6084# m1_n5428_n5842# pfet$272
Xpfet$275_19 vdd vdd m1_n3884_n9085# m1_n5427_n8573# pfet$275
Xpfet$272_3 vdd vdd m1_n5868_n3849# fref pfet$272
Xpfet$270_0 vdd vdd m1_5464_n5483# m1_5895_n8089# pfet$270
Xnfet$296_0 m1_n3884_n11124# vss m1_n3098_n10720# vss nfet$296
Xpfet$270_1 vdd vdd m1_4978_n5483# m1_5464_n5483# pfet$270
Xnfet$296_1 m1_n3884_n9085# vss m1_n3098_n9135# vss nfet$296
Xnfet$289_0 m1_5895_n8089# vss m1_5464_n5483# vss nfet$289
Xnfet$289_1 m1_5464_n5483# vss m1_4978_n5483# vss nfet$289
Xnfet$294_0 m1_2556_n10129# m1_2556_n10129# vss vss m1_3015_n10205# vss nfet$294
Xnfet$294_1 m1_1452_n8889# m1_1452_n8889# m1_1096_n9089# m1_1096_n9089# m1_1550_n9245#
+ vss nfet$294
Xnfet$287_0 m1_2779_n3533# vss up vss nfet$287
Xnfet$294_2 m1_2068_n8889# m1_2068_n8889# vss vss m1_1550_n9245# vss nfet$294
Xnfet$287_1 m1_2779_n3533# vss m1_3349_n5165# vss nfet$287
Xnfet$287_2 m1_2758_n8889# vss m1_2068_n5361# vss nfet$287
Xnfet$294_3 m1_2068_n8889# m1_2068_n8889# m1_2779_n10883# m1_2779_n10883# m1_3015_n10205#
+ vss nfet$294
Xpfet$277_0 m1_n4677_n8889# vdd vdd m1_n1925_n10720# pfet$277
Xnfet$292_0 m1_n4678_n3849# m1_n4678_n3849# m1_n5428_n3533# m1_n5428_n3533# m1_n5192_n4205#
+ vss nfet$292
Xnfet$287_3 m1_832_n5785# vss m1_1452_n5483# vss nfet$287
Xnfet$285_0 m1_n3885_n4045# m1_832_n5785# m1_1096_n5165# vss nfet$285
Xnfet$294_4 m1_n4677_n10522# m1_n4677_n10522# m1_n5427_n10882# m1_n5427_n10882# m1_n5191_n10204#
+ vss nfet$294
Xnfet$292_1 m1_n5650_n4045# m1_n5650_n4045# vss vss m1_n5192_n4205# vss nfet$292
Xpfet$277_1 m1_n1925_n10720# vdd vdd m1_n3098_n10720# pfet$277
Xnfet$287_4 vdd vss m1_1095_n4045# vss nfet$287
Xnfet$294_5 m1_n5649_n11124# m1_n5649_n11124# vss vss m1_n5191_n10204# vss nfet$294
Xnfet$285_1 m1_n3885_n4045# m1_1452_n5483# m1_2556_n4049# vss nfet$285
Xpfet$277_2 m1_n4677_n10522# vdd vdd m1_n1925_n9135# pfet$277
Xnfet$292_2 m1_n4678_n5482# m1_n4678_n5482# m1_n5428_n5842# m1_n5428_n5842# m1_n5192_n5164#
+ vss nfet$292
Xnfet$285_2 m1_n3885_n6084# m1_1095_n4045# m1_832_n5785# vss nfet$285
Xnfet$294_6 m1_n4677_n8889# m1_n4677_n8889# m1_n5427_n8573# m1_n5427_n8573# m1_n5191_n9245#
+ vss nfet$294
Xnfet$292_3 m1_n5868_n3849# m1_n5868_n3849# vss vss m1_n5192_n5164# vss nfet$292
Xpfet$275_0 vdd vdd m1_2779_n10883# m1_2068_n8889# pfet$275
Xpfet$277_3 m1_n1925_n9135# vdd vdd m1_n3098_n9135# pfet$277
Xnfet$290_0 m1_n1926_n4095# m1_n3099_n4095# vss vss nfet$290
Xnfet$294_7 m1_n5867_n10544# m1_n5867_n10544# vss vss m1_n5191_n9245# vss nfet$294
Xnfet$285_3 m1_n3885_n6084# m1_2556_n4049# m1_3349_n5165# vss nfet$285
Xpfet$275_1 vdd m1_2779_n10883# vdd m1_2556_n10129# pfet$275
Xnfet$290_1 m1_n4678_n3849# m1_n1926_n5680# vss vss nfet$290
Xpfet$268_0 vdd vdd m1_3349_n5165# m1_2779_n3533# pfet$268
Xpfet$275_2 vdd m1_1095_n11125# m1_832_n8573# m1_n3884_n11124# pfet$275
Xnfet$290_2 m1_n1926_n5680# m1_n3099_n5680# vss vss nfet$290
Xpfet$268_1 vdd vdd up m1_2779_n3533# pfet$268
Xpfet$268_2 vdd vdd m1_2068_n5361# m1_2758_n8889# pfet$268
Xpfet$275_3 vdd m1_1452_n8889# m1_2556_n10129# m1_n3884_n9085# pfet$275
Xnfet$290_3 m1_n4678_n5482# m1_n1926_n4095# vss vss nfet$290
Xpfet$273_0 vdd m1_n5428_n3533# vdd m1_n5650_n4045# pfet$273
Xpfet$275_4 vdd vdd m1_1452_n8889# m1_832_n8573# pfet$275
Xpfet$268_3 vdd vdd m1_1452_n5483# m1_832_n5785# pfet$268
Xpfet$266_0 vdd m1_832_n5785# m1_1096_n5165# m1_n3885_n6084# pfet$266
Xpfet$273_1 vdd vdd m1_n5428_n3533# m1_n4678_n3849# pfet$273
Xpfet$268_4 vdd vdd m1_1095_n4045# vdd pfet$268
Xpfet$275_5 vdd vdd m1_1095_n11125# vdd pfet$275
Xpfet$266_1 vdd m1_1452_n5483# m1_2556_n4049# m1_n3885_n6084# pfet$266
Xpfet$273_2 vdd m1_n5428_n5842# vdd m1_n5868_n3849# pfet$273
Xpfet$266_2 vdd m1_1095_n4045# m1_832_n5785# m1_n3885_n4045# pfet$266
Xpfet$275_6 vdd vdd m1_1096_n9089# m1_1452_n8889# pfet$275
Xpfet$273_3 vdd vdd m1_n5428_n5842# m1_n4678_n5482# pfet$273
Xpfet$271_0 m1_n1926_n4095# vdd vdd m1_n3099_n4095# pfet$271
Xnfet$297_0 m1_n4677_n8889# m1_n1925_n10720# vss vss nfet$297
Xpfet$275_7 vdd m1_832_n8573# m1_1096_n9089# m1_n3884_n9085# pfet$275
Xpfet$266_3 vdd m1_2556_n4049# m1_3349_n5165# m1_n3885_n4045# pfet$266
Xpfet$271_1 m1_n4678_n3849# vdd vdd m1_n1926_n5680# pfet$271
Xnfet$297_1 m1_n1925_n10720# m1_n3098_n10720# vss vss nfet$297
Xpfet$275_8 vdd m1_1096_n9089# vdd m1_2068_n8889# pfet$275
Xpfet$271_2 m1_n1926_n5680# vdd vdd m1_n3099_n5680# pfet$271
Xpfet$275_9 vdd vdd m1_2068_n8889# m1_2758_n8889# pfet$275
Xnfet$297_2 m1_n4677_n10522# m1_n1925_n9135# vss vss nfet$297
Xpfet$271_3 m1_n4678_n5482# vdd vdd m1_n1926_n4095# pfet$271
Xnfet$297_3 m1_n1925_n9135# m1_n3098_n9135# vss vss nfet$297
Xnfet$295_0 m1_n3884_n9085# m1_1095_n11125# m1_832_n8573# vss nfet$295
Xnfet$295_1 m1_n3884_n11124# m1_1452_n8889# m1_2556_n10129# vss nfet$295
Xnfet$288_0 m1_4978_n5483# vss m1_2758_n8889# vss nfet$288
Xnfet$295_10 m1_n5867_n10544# vss m1_n5649_n11124# vss nfet$295
Xnfet$295_2 m1_832_n8573# vss m1_1452_n8889# vss nfet$295
Xnfet$295_11 fdiv vss m1_n5867_n10544# vss nfet$295
Xnfet$295_3 vdd vss m1_1095_n11125# vss nfet$295
Xpfet$278_0 vdd m1_5895_n8089# vdd down pfet$278
Xnfet$295_12 m1_n5427_n8573# vss m1_n3884_n9085# vss nfet$295
Xnfet$293_0 m1_n3885_n4045# vss m1_n3099_n4095# vss nfet$293
Xnfet$295_4 m1_n3884_n11124# m1_832_n8573# m1_1096_n9089# vss nfet$295
Xnfet$286_0 m1_2068_n5361# m1_2068_n5361# vss vss m1_1550_n5165# vss nfet$286
Xpfet$278_1 vdd vdd m1_5895_n8089# up pfet$278
Xnfet$293_1 m1_n3885_n6084# vss m1_n3099_n5680# vss nfet$293
Xpfet$275_20 vdd m1_n5427_n8573# vdd m1_n5867_n10544# pfet$275
Xnfet$286_1 m1_1452_n5483# m1_1452_n5483# m1_1096_n5165# m1_1096_n5165# m1_1550_n5165#
+ vss nfet$286
Xnfet$295_5 m1_2758_n8889# vss m1_2068_n8889# vss nfet$295
Xnfet$295_6 m1_2779_n10883# vss down vss nfet$295
Xpfet$275_10 vdd vdd m1_3349_n9089# m1_2779_n10883# pfet$275
Xnfet$286_2 m1_2556_n4049# m1_2556_n4049# vss vss m1_3015_n4205# vss nfet$286
Xnfet$291_0 m1_n5428_n3533# vss m1_n3885_n4045# vss nfet$291
Xpfet$276_0 vdd vdd m1_n3098_n10720# m1_n3884_n11124# pfet$276
Xpfet$275_11 vdd vdd down m1_2779_n10883# pfet$275
Xnfet$286_3 m1_2068_n5361# m1_2068_n5361# m1_2779_n3533# m1_2779_n3533# m1_3015_n4205#
+ vss nfet$286
Xnfet$295_7 m1_2779_n10883# vss m1_3349_n9089# vss nfet$295
Xpfet$276_1 vdd vdd m1_n3098_n9135# m1_n3884_n9085# pfet$276
Xnfet$291_1 m1_n5868_n3849# vss m1_n5650_n4045# vss nfet$291
Xpfet$269_0 vdd vdd m1_2758_n8889# m1_4978_n5483# pfet$269
Xnfet$295_8 m1_n3884_n9085# m1_2556_n10129# m1_3349_n9089# vss nfet$295
Xpfet$275_12 vdd m1_2556_n10129# m1_3349_n9089# m1_n3884_n11124# pfet$275
Xnfet$291_2 m1_n5428_n5842# vss m1_n3885_n6084# vss nfet$291
Xpfet$275_13 vdd vdd m1_n5427_n8573# m1_n4677_n8889# pfet$275
Xnfet$295_9 m1_n5427_n10882# vss m1_n3884_n11124# vss nfet$295
Xnfet$291_3 fref vss m1_n5868_n3849# vss nfet$291
Xpfet$274_0 vdd vdd m1_n3099_n4095# m1_n3885_n4045# pfet$274
Xpfet$275_14 vdd vdd m1_n3884_n11124# m1_n5427_n10882# pfet$275
Xpfet$274_1 vdd vdd m1_n3099_n5680# m1_n3885_n6084# pfet$274
Xpfet$267_0 vdd vdd m1_1096_n5165# m1_1452_n5483# pfet$267
Xpfet$275_15 vdd m1_n5427_n10882# vdd m1_n5649_n11124# pfet$275
Xpfet$267_1 vdd m1_1096_n5165# vdd m1_2068_n5361# pfet$267
Xpfet$275_16 vdd vdd m1_n5427_n10882# m1_n4677_n10522# pfet$275
Xpfet$267_2 vdd m1_2779_n3533# vdd m1_2556_n4049# pfet$267
Xpfet$272_0 vdd vdd m1_n3885_n4045# m1_n5428_n3533# pfet$272
.ends

.subckt pfet$279 a_254_0# a_348_560# w_n180_n88# a_414_0# a_n92_0# a_94_0# a_574_0#
+ a_508_560# a_188_560# a_28_560#
X0 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$299 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt BIAS vdd vss res 200p1 200p2 100n 200n
Xpfet$279_10 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$279
Xpfet$279_11 vdd res vdd 200n vdd 200n vdd res res res pfet$279
Xpfet$279_1 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$279
Xpfet$279_0 vdd res vdd 200n vdd 200n vdd res res res pfet$279
Xpfet$279_13 vdd res vdd res vdd res vdd res res res pfet$279
Xpfet$279_12 vdd res vdd 100n vdd 100n vdd res res res pfet$279
Xpfet$279_2 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$279
Xpfet$279_14 vdd res vdd 200n vdd 200n vdd res res res pfet$279
Xpfet$279_3 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$279
Xpfet$279_15 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$279
Xpfet$279_4 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$279
Xpfet$279_5 vdd res vdd 200n vdd 200n vdd res res res pfet$279
Xpfet$279_6 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$279
Xpfet$279_7 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$279
Xpfet$279_8 vdd res vdd res vdd res vdd res res res pfet$279
Xpfet$279_9 vdd res vdd 100n vdd 100n vdd res res res pfet$279
Xnfet$299_0 m1_27_n1423# vss 200p1 m1_27_n1423# vss 200p1 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$299
Xnfet$299_1 vss vss vss vss vss vss vss vss vss vss nfet$299
Xnfet$299_2 m1_27_n1423# vss 200p2 m1_27_n1423# vss 200p2 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$299
Xnfet$299_3 vss vss vss vss vss vss vss vss vss vss nfet$299
Xnfet$299_4 m1_27_n1423# vss 200p2 m1_27_n1423# vss 200p2 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$299
Xnfet$299_5 m1_27_n1423# vss 200p1 m1_27_n1423# vss 200p1 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$299
Xnfet$299_6 m1_27_n1423# vss m1_27_n1423# m1_27_n1423# vss m1_27_n1423# m1_27_n1423#
+ vss m1_27_n1423# vss nfet$299
Xnfet$299_7 m1_27_n1423# vss m1_27_n1423# m1_27_n1423# vss m1_27_n1423# m1_27_n1423#
+ vss m1_27_n1423# vss nfet$299
.ends

.subckt nfet$300 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.5u
.ends

.subckt cap_mim m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
.ends

.subckt pfet$282 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$280 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=9.75p pd=31.3u as=9.75p ps=31.3u w=15u l=0.5u
.ends

.subckt nfet$301 a_n84_0# a_38_n132# a_138_0# VSUBS
X0 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.5u
.ends

.subckt pfet$281 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=9.75p pd=31.3u as=9.75p ps=31.3u w=15u l=0.5u
.ends

.subckt nfet$302 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt CSRVCO_20250823 vctrl vosc vdd vss
Xnfet$300_0 m1_n9838_266# m1_n12754_674# m1_n9352_266# vss nfet$300
Xnfet$300_1 vctrl vss m1_n12268_985# vss nfet$300
Xnfet$300_2 vctrl vss m1_n14283_186# vss nfet$300
Xnfet$300_3 vctrl vss m1_n13794_186# vss nfet$300
Xnfet$300_4 vctrl vss m1_n13240_368# vss nfet$300
Xnfet$300_5 vctrl vss m1_n12754_674# vss nfet$300
Xnfet$300_6 vctrl m1_n16019_266# vss vss nfet$300
Xnfet$300_7 vctrl vss m1_n15245_186# vss nfet$300
Xnfet$300_8 vctrl vss m1_n14765_186# vss nfet$300
Xnfet$300_9 m1_n10324_266# m1_n13240_368# m1_n9838_266# vss nfet$300
Xcap_mim_0 vss m1_n11296_266# cap_mim
Xcap_mim_1 vss m1_n10810_266# cap_mim
Xpfet$282_0 vdd vdd vosc m1_n8380_274# pfet$282
Xcap_mim_2 vss m1_n10324_266# cap_mim
Xpfet$282_1 vdd vdd m1_n8380_274# m1_n11916_1270# pfet$282
Xcap_mim_3 vss m1_n11916_1270# cap_mim
Xcap_mim_5 vss m1_n9838_266# cap_mim
Xcap_mim_4 vss m1_n9352_266# cap_mim
Xpfet$280_0 vdd vdd m1_n12264_2422# m1_n16019_266# pfet$280
Xnfet$300_10 m1_n9352_266# m1_n12268_985# m1_n11916_1270# vss nfet$300
Xcap_mim_6 vss m1_n11782_266# cap_mim
Xpfet$280_1 vdd vdd m1_n14208_3657# m1_n16019_266# pfet$280
Xnfet$300_11 m1_n11916_1270# m1_n15245_186# m1_n11782_266# vss nfet$300
Xnfet$301_0 vss vss vss vss nfet$301
Xpfet$280_2 vdd vdd m1_n13722_3340# m1_n16019_266# pfet$280
Xnfet$301_1 vss vss vss vss nfet$301
Xnfet$300_12 m1_n11782_266# m1_n14765_186# m1_n11296_266# vss nfet$300
Xpfet$280_3 vdd m1_n16019_266# vdd m1_n16019_266# pfet$280
Xnfet$300_13 m1_n11296_266# m1_n14283_186# m1_n10810_266# vss nfet$300
Xpfet$280_4 vdd vdd m1_n13236_3035# m1_n16019_266# pfet$280
Xnfet$300_14 m1_n10810_266# m1_n13794_186# m1_n10324_266# vss nfet$300
Xpfet$280_6 vdd vdd m1_n12750_2729# m1_n16019_266# pfet$280
Xpfet$280_5 vdd vdd m1_n14693_3963# m1_n16019_266# pfet$280
Xpfet$280_7 vdd vdd m1_n15180_4275# m1_n16019_266# pfet$280
Xpfet$280_8 vdd m1_n13236_3035# m1_n9838_266# m1_n10324_266# pfet$280
Xpfet$280_9 vdd m1_n12750_2729# m1_n9352_266# m1_n9838_266# pfet$280
Xpfet$280_10 vdd m1_n14208_3657# m1_n10810_266# m1_n11296_266# pfet$280
Xpfet$280_11 vdd m1_n12264_2422# m1_n11916_1270# m1_n9352_266# pfet$280
Xpfet$280_12 vdd m1_n14693_3963# m1_n11296_266# m1_n11782_266# pfet$280
Xpfet$280_13 vdd m1_n13722_3340# m1_n10324_266# m1_n10810_266# pfet$280
Xpfet$281_0 vdd vdd vdd vdd pfet$281
Xpfet$281_1 vdd vdd vdd vdd pfet$281
Xpfet$280_14 vdd m1_n15180_4275# m1_n11782_266# m1_n11916_1270# pfet$280
Xnfet$302_0 m1_n8380_274# vss vosc vss nfet$302
Xnfet$302_1 m1_n11916_1270# vss m1_n8380_274# vss nfet$302
.ends

.subckt asc_hysteresis_buffer$6 vss in vdd out
Xpfet$235_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd
+ m1_884_42# m1_884_42# pfet$235
Xnfet$257_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$257
Xnfet$255_0 m1_348_648# vss m1_884_42# vss nfet$255
Xpfet$238_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$238
Xpfet$236_0 vdd vdd m1_884_42# m1_348_648# pfet$236
Xnfet$258_0 m1_1156_42# vss m1_884_42# vss nfet$258
Xnfet$256_0 in vss m1_348_648# vss nfet$256
Xnfet$254_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$254
Xpfet$239_0 vdd vdd m1_884_42# m1_1156_42# pfet$239
Xpfet$237_0 vdd vdd m1_348_648# in pfet$237
.ends

.subckt top_level_20250912_nosc i_cp_100u div_def div_prc_s8 div_prc_s7 div_prc_s6
+ div_prc_s5 div_prc_s4 div_prc_s3 div_prc_s2 div_prc_s1 div_prc_s0 div_in div_swc_s0
+ div_swc_s1 div_swc_s2 div_swc_s3 div_swc_s4 div_swc_s5 div_swc_s6 div_swc_s7 div_swc_s8
+ lock ref ext_pfd_div ext_pfd_ref ext_pfd_up ext_pfd_down mx_pfd_s1 mx_pfd_s0 down
+ cp_s1 cp_s2 cp_s3 cp_s4 filter_in out filter_out mx_vco_s0 mx_vco_s1 div_rpc_s0
+ div_rsc_s0 div_rsc_s1 div_rpc_s1 div_rsc_s2 div_rpc_s2 div_rsc_s3 div_rsc_s4 div_rsc_s5
+ div_rsc_s6 div_rsc_s7 div_rsc_s8 div_rpc_s3 div_rpc_s4 div_rpc_s5 div_rpc_s6 div_rpc_s7
+ div_rpc_s8 mx_ref_s1 mx_ref_s0 up ext_vco_out vdd vss ext_vco_in div_out
Xasc_drive_buffer_up_0 vss asc_drive_buffer_up_0/out xp_3_1_MUX_2/OUT_1 vdd asc_drive_buffer_up
Xasc_dual_psd_def_20250809_0 vdd vss div_prc_s0 div_prc_s1 div_prc_s2 div_prc_s3 div_prc_s4
+ div_prc_s5 div_prc_s6 div_prc_s7 div_prc_s8 xp_3_1_MUX_4/OUT_1 div_swc_s0 div_swc_s1
+ div_swc_s2 div_swc_s3 div_swc_s4 div_swc_s5 div_swc_s6 div_swc_s7 div_swc_s8 asc_drive_buffer_0/in
+ div_def asc_dual_psd_def_20250809
Xasc_drive_buffer_0 vss asc_drive_buffer_0/in vdd div_in asc_drive_buffer
Xasc_drive_buffer_1 vss xp_3_1_MUX_0/OUT_1 vdd out asc_drive_buffer
Xasc_drive_buffer_2 vss xp_3_1_MUX_4/OUT_1 vdd div_out asc_drive_buffer
Xasc_drive_buffer_3 vss asc_drive_buffer_3/in vdd lock asc_drive_buffer
Xasc_lock_detector_20250826_0 xp_3_1_MUX_3/OUT_1 vdd xp_3_1_MUX_4/OUT_1 asc_drive_buffer_3/in
+ vss asc_lock_detector_20250826
Xasc_drive_buffer_4 vss xp_3_1_MUX_2/OUT_1 vdd up asc_drive_buffer
Xasc_drive_buffer_5 vss xp_3_1_MUX_5/OUT_1 vdd down asc_drive_buffer
Xasc_drive_buffer_6 vss xp_3_1_MUX_5/OUT_1 vdd asc_drive_buffer_6/out asc_drive_buffer
Xxp_3_1_MUX_0 mx_vco_s0 mx_vco_s1 vdd vss xp_3_1_MUX_0/OUT_1 xp_3_1_MUX_0/C_1 xp_3_1_MUX_0/B_1
+ ext_vco_out xp_3_1_MUX
Xxp_3_1_MUX_1 mx_vco_s0 mx_vco_s1 vdd vss filter_out xp_3_1_MUX_1/C_1 xp_3_1_MUX_1/B_1
+ ext_vco_in xp_3_1_MUX
Xxp_3_1_MUX_2 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX_2/OUT_1 xp_3_1_MUX_2/C_1 xp_3_1_MUX_2/B_1
+ ext_pfd_up xp_3_1_MUX
Xxp_3_1_MUX_3 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX_3/OUT_1 xp_3_1_MUX_3/C_1 xp_3_1_MUX_3/B_1
+ ext_pfd_ref xp_3_1_MUX
Xxp_3_1_MUX_4 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX_4/OUT_1 xp_3_1_MUX_4/C_1 xp_3_1_MUX_4/B_1
+ ext_pfd_div xp_3_1_MUX
Xxp_programmable_basic_pump_0 asc_drive_buffer_up_0/out vdd cp_s1 cp_s2 cp_s3 cp_s4
+ asc_drive_buffer_6/out filter_in BIAS_0/100n vss xp_programmable_basic_pump
Xasc_hysteresis_buffer$5_0 vss xp_3_1_MUX$4_1/OUT_1 vdd xp_3_1_MUX_3/OUT_1 asc_hysteresis_buffer$5
Xxp_3_1_MUX_5 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX_5/OUT_1 xp_3_1_MUX_5/C_1 xp_3_1_MUX_5/B_1
+ ext_pfd_down xp_3_1_MUX
Xxp_3_1_MUX$4_0 mx_ref_s0 mx_ref_s1 vdd vss xp_3_1_MUX$4_0/OUT_1 xp_3_1_MUX$4_1/C_1
+ xp_3_1_MUX$4_0/B_1 xp_3_1_MUX$4_0/A_1 xp_3_1_MUX$4
Xxp_3_1_MUX$4_1 mx_ref_s0 mx_ref_s1 vdd vss xp_3_1_MUX$4_1/OUT_1 xp_3_1_MUX$4_1/C_1
+ xp_3_1_MUX$4_1/B_1 xp_3_1_MUX$4_1/A_1 xp_3_1_MUX$4
Xasc_dual_psd_def_20250809$4_0 vdd vss div_rpc_s0 div_rpc_s1 div_rpc_s2 div_rpc_s3
+ div_rpc_s4 div_rpc_s5 div_rpc_s6 div_rpc_s7 div_rpc_s8 xp_3_1_MUX$4_1/B_1 div_rsc_s0
+ div_rsc_s1 div_rsc_s2 div_rsc_s3 div_rsc_s4 div_rsc_s5 div_rsc_s6 div_rsc_s7 div_rsc_s8
+ xp_3_1_MUX$4_0/B_1 vss asc_dual_psd_def_20250809$4
Xasc_drive_buffer$4_0 vss xp_3_1_MUX_0/OUT_1 vdd asc_drive_buffer_0/in asc_drive_buffer$4
Xasc_PFD_DFF_20250831_0 vss xp_3_1_MUX_3/C_1 xp_3_1_MUX_5/C_1 xp_3_1_MUX_2/C_1 vdd
+ xp_3_1_MUX_4/C_1 asc_PFD_DFF_20250831
XBIAS_0 vdd vss i_cp_100u BIAS_0/200p1 BIAS_0/200p2 BIAS_0/100n BIAS_0/200n BIAS
Xasc_PFD_DFF_20250831_1 vss xp_3_1_MUX_3/B_1 xp_3_1_MUX_2/B_1 xp_3_1_MUX_5/B_1 vdd
+ xp_3_1_MUX_4/B_1 asc_PFD_DFF_20250831
XCSRVCO_20250823_0 xp_3_1_MUX_1/C_1 xp_3_1_MUX_0/C_1 vdd vss CSRVCO_20250823
Xasc_hysteresis_buffer$6_0 vss ref vdd xp_3_1_MUX$4_0/OUT_1 asc_hysteresis_buffer$6
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__and2_1 A1 A2 VDD VSS Z VNW VPW
X0 VDD A2 a_36_201# VNW pfet_05v0 ad=0.5054p pd=2.57u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1 a_244_201# A1 a_36_201# VPW nfet_05v0 ad=0.1056p pd=0.98u as=0.2904p ps=2.2u w=0.66u l=0.6u
X2 Z a_36_201# VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.3894p ps=2.06u w=1.32u l=0.6u
X3 Z a_36_201# VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.5054p ps=2.57u w=1.83u l=0.5u
X4 VSS A2 a_244_201# VPW nfet_05v0 ad=0.3894p pd=2.06u as=0.1056p ps=0.98u w=0.66u l=0.6u
X5 a_36_201# A1 VDD VNW pfet_05v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__latq_1 D E Q VDD VSS VNW VPW
X0 VSS a_1020_652# Q VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X1 a_504_110# a_36_92# VDD VNW pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X2 VDD a_1020_652# Q VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X3 a_1264_107# a_36_92# a_1020_652# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X4 VSS E a_36_92# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X5 VSS a_1364_532# a_1264_107# VPW nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X6 VDD E a_36_92# VNW pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X7 VDD a_1364_532# a_1224_652# VNW pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X8 a_872_652# D VDD VNW pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X9 a_1364_532# a_1020_652# VDD VNW pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X10 a_1020_652# a_504_110# a_872_107# VPW nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X11 a_872_107# D VSS VPW nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X12 a_1020_652# a_36_92# a_872_652# VNW pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X13 a_504_110# a_36_92# VSS VPW nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X14 a_1364_532# a_1020_652# VSS VPW nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X15 a_1224_652# a_504_110# a_1020_652# VNW pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt DFF_2phase_1 VDDd D PHI_2 PHI_1 Q VSSd
Xgf180mcu_fd_sc_mcu9t5v0__latq_1_0 gf180mcu_fd_sc_mcu9t5v0__latq_1_1/Q PHI_2 Q VDDd
+ VSSd VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1
Xgf180mcu_fd_sc_mcu9t5v0__latq_1_1 D PHI_1 gf180mcu_fd_sc_mcu9t5v0__latq_1_1/Q VDDd
+ VSSd VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1 I VDD VSS ZN VNW VPW
X0 ZN I VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__or2_1 A1 A2 VDD VSS Z VNW VPW
X0 a_255_756# A1 a_67_756# VNW pfet_05v0 ad=0.2379p pd=1.435u as=0.4026p ps=2.71u w=0.915u l=0.5u
X1 VSS A2 a_67_756# VPW nfet_05v0 ad=0.3828p pd=2.08u as=0.1716p ps=1.18u w=0.66u l=0.6u
X2 VDD A2 a_255_756# VNW pfet_05v0 ad=0.57645p pd=2.69u as=0.2379p ps=1.435u w=0.915u l=0.5u
X3 Z a_67_756# VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.3828p ps=2.08u w=1.32u l=0.6u
X4 Z a_67_756# VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.57645p ps=2.69u w=1.83u l=0.5u
X5 a_67_756# A1 VSS VPW nfet_05v0 ad=0.1716p pd=1.18u as=0.2904p ps=2.2u w=0.66u l=0.6u
.ends

.subckt Register_unitcell out default d en phi2 q phi1 VSSd VDDd
Xgf180mcu_fd_sc_mcu9t5v0__and2_1_1 q en VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1_0/A2
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1
XDFF_2phase_1_0 VDDd d phi2 phi1 q VSSd DFF_2phase_1
Xgf180mcu_fd_sc_mcu9t5v0__inv_1_0 en VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1_0/ZN
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
Xgf180mcu_fd_sc_mcu9t5v0__or2_1_0 gf180mcu_fd_sc_mcu9t5v0__or2_1_0/A1 gf180mcu_fd_sc_mcu9t5v0__or2_1_0/A2
+ VDDd VSSd out VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1
Xgf180mcu_fd_sc_mcu9t5v0__and2_1_0 gf180mcu_fd_sc_mcu9t5v0__inv_1_0/ZN default VDDd
+ VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1_0/A1 VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1
.ends

.subckt SRegister_10 out[1] out[2] out[3] out[9] default10 default9 default8 default7
+ default6 default5 default4 default3 default2 default1 d q out[6] out[4] out[10]
+ out[7] out[5] phi2 out[8] VDDd en VSSd phi1
XRegister_unitcell_0 out[2] default2 Register_unitcell_6/q en phi2 Register_unitcell_7/d
+ phi1 VSSd VDDd Register_unitcell
XRegister_unitcell_1 out[6] default6 Register_unitcell_9/q en phi2 Register_unitcell_2/d
+ phi1 VSSd VDDd Register_unitcell
XRegister_unitcell_2 out[7] default7 Register_unitcell_2/d en phi2 Register_unitcell_3/d
+ phi1 VSSd VDDd Register_unitcell
XRegister_unitcell_3 out[8] default8 Register_unitcell_3/d en phi2 Register_unitcell_4/d
+ phi1 VSSd VDDd Register_unitcell
XRegister_unitcell_5 out[10] default10 Register_unitcell_5/d en phi2 q phi1 VSSd VDDd
+ Register_unitcell
XRegister_unitcell_4 out[9] default9 Register_unitcell_4/d en phi2 Register_unitcell_5/d
+ phi1 VSSd VDDd Register_unitcell
XRegister_unitcell_6 out[1] default1 d en phi2 Register_unitcell_6/q phi1 VSSd VDDd
+ Register_unitcell
XRegister_unitcell_7 out[3] default3 Register_unitcell_7/d en phi2 Register_unitcell_8/d
+ phi1 VSSd VDDd Register_unitcell
XRegister_unitcell_8 out[4] default4 Register_unitcell_8/d en phi2 Register_unitcell_9/d
+ phi1 VSSd VDDd Register_unitcell
XRegister_unitcell_9 out[5] default5 Register_unitcell_9/d en phi2 Register_unitcell_9/q
+ phi1 VSSd VDDd Register_unitcell
.ends

.subckt pfet$192 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt nfet$208 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt pfet$195 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$209 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$193 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt nfet$207 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt nfet$210 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$194 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt qw_NOLclk CLK VDDd VSSd PHI_1 PHI_2
Xpfet$192_1 VDDd VDDd m1_13930_1818# PHI_2 pfet$192
Xnfet$208_2 m1_12351_431# m1_15103_1818# VSSd VSSd nfet$208
Xnfet$208_3 m1_15103_1818# m1_13930_1818# VSSd VSSd nfet$208
Xpfet$195_0 VDDd m1_11601_71# VDDd m1_11379_n171# pfet$195
Xpfet$195_1 VDDd VDDd m1_11601_71# m1_12351_431# pfet$195
Xpfet$195_3 VDDd VDDd m1_11601_2380# m1_12351_2064# pfet$195
Xpfet$195_2 VDDd m1_11601_2380# VDDd m1_11161_409# pfet$195
Xnfet$209_0 m1_11601_71# VSSd PHI_1 VSSd nfet$209
Xnfet$209_2 m1_11601_2380# VSSd PHI_2 VSSd nfet$209
Xnfet$209_1 m1_11161_409# VSSd m1_11379_n171# VSSd nfet$209
Xpfet$193_0 m1_12351_2064# VDDd VDDd m1_15103_233# pfet$193
Xpfet$193_1 m1_15103_233# VDDd VDDd m1_13930_233# pfet$193
Xpfet$193_2 m1_12351_431# VDDd VDDd m1_15103_1818# pfet$193
Xnfet$209_3 CLK VSSd m1_11161_409# VSSd nfet$209
Xnfet$207_0 PHI_1 VSSd m1_13930_233# VSSd nfet$207
Xpfet$193_3 m1_15103_1818# VDDd VDDd m1_13930_1818# pfet$193
Xnfet$207_1 PHI_2 VSSd m1_13930_1818# VSSd nfet$207
Xnfet$210_0 m1_12351_431# m1_12351_431# m1_11601_71# m1_11601_71# m1_11837_749# VSSd
+ nfet$210
Xnfet$210_1 m1_11379_n171# m1_11379_n171# VSSd VSSd m1_11837_749# VSSd nfet$210
Xnfet$210_2 m1_12351_2064# m1_12351_2064# m1_11601_2380# m1_11601_2380# m1_11837_1708#
+ VSSd nfet$210
Xnfet$210_3 m1_11161_409# m1_11161_409# VSSd VSSd m1_11837_1708# VSSd nfet$210
Xpfet$194_0 VDDd VDDd PHI_1 m1_11601_71# pfet$194
Xpfet$194_1 VDDd VDDd m1_11379_n171# m1_11161_409# pfet$194
Xpfet$194_2 VDDd VDDd PHI_2 m1_11601_2380# pfet$194
Xnfet$208_0 m1_12351_2064# m1_15103_233# VSSd VSSd nfet$208
Xpfet$194_3 VDDd VDDd m1_11161_409# CLK pfet$194
Xnfet$208_1 m1_15103_233# m1_13930_233# VSSd VSSd nfet$208
Xpfet$192_0 VDDd VDDd m1_13930_233# PHI_1 pfet$192
.ends

.subckt pfet a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$204 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$202 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$188 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$186 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0#
+ a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$203 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$201 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$189 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$187 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt asc_hysteresis_buffer vss in vdd out
Xpfet_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd m1_884_42#
+ m1_884_42# pfet
Xnfet$204_0 m1_1156_42# vss m1_884_42# vss nfet$204
Xnfet$202_0 in vss m1_348_648# vss nfet$202
Xpfet$188_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$188
Xpfet$186_0 vdd vdd m1_884_42# m1_348_648# pfet$186
Xnfet_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42# vss
+ m1_884_42# vss nfet
Xnfet$203_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$203
Xnfet$201_0 m1_348_648# vss m1_884_42# vss nfet$201
Xpfet$189_0 vdd vdd m1_884_42# m1_1156_42# pfet$189
Xpfet$187_0 vdd vdd m1_348_648# in pfet$187
.ends

.subckt nfet$206 a_30_n132# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$190 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=2.6p pd=9.3u as=2.6p ps=9.3u w=4u l=0.28u
.ends

.subckt pfet$191 a_28_460# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_460# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt nfet$205 a_n84_0# a_94_0# a_30_460# VSUBS
X0 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt SCHMITT VDD VSS IN OUT
Xnfet$206_0 OUT m1_592_402# VDD VSS nfet$206
Xpfet$190_0 IN VDD m1_596_1544# OUT pfet$190
Xpfet$190_1 IN VDD VDD m1_596_1544# pfet$190
Xpfet$191_0 OUT VDD m1_596_1544# VSS pfet$191
Xnfet$205_0 m1_592_402# OUT IN VSS nfet$205
Xnfet$205_1 VSS m1_592_402# IN VSS nfet$205
.ends

.subckt scan_chain VDDd ENd DATAd CLKd out[1] out[2] out[3] out[4] out[5] out[6] out[7]
+ out[8] out[9] out[10] out[20] out[19] out[18] out[17] out[16] out[15] out[14] out[13]
+ out[12] out[11] out[21] out[22] out[23] out[24] out[25] out[26] out[27] out[28]
+ out[29] out[30] out[40] out[39] out[38] out[37] out[36] out[35] out[34] out[33]
+ out[32] out[31] out[41] out[42] out[43] out[44] out[45] out[46] out[47] out[48]
+ out[49] out[50] VSSd
XSRegister_10_1 out[11] out[12] out[13] out[19] VSSd VSSd VSSd VSSd VSSd VSSd VSSd
+ VSSd VSSd VSSd SRegister_10_4/q SRegister_10_3/d out[16] out[14] out[20] out[17]
+ out[15] qw_NOLclk_0/PHI_2 out[18] VDDd SRegister_10_4/en VSSd qw_NOLclk_0/PHI_1
+ SRegister_10
XSRegister_10_2 out[41] out[42] out[43] out[49] VSSd VSSd VSSd VSSd VDDd VSSd VSSd
+ VDDd VDDd VSSd SRegister_10_2/d SRegister_10_2/q out[46] out[44] out[50] out[47]
+ out[45] qw_NOLclk_0/PHI_2 out[48] VDDd SRegister_10_4/en VSSd qw_NOLclk_0/PHI_1
+ SRegister_10
Xqw_NOLclk_0 SCHMITT_0/OUT VDDd VSSd qw_NOLclk_0/PHI_1 qw_NOLclk_0/PHI_2 qw_NOLclk
XSRegister_10_3 out[21] out[22] out[23] out[29] VSSd VSSd VSSd VSSd VSSd VSSd VSSd
+ VSSd VSSd VSSd SRegister_10_3/d SRegister_10_3/q out[26] out[24] out[30] out[27]
+ out[25] qw_NOLclk_0/PHI_2 out[28] VDDd SRegister_10_4/en VSSd qw_NOLclk_0/PHI_1
+ SRegister_10
XSRegister_10_4 out[1] out[2] out[3] out[9] VSSd VSSd VSSd VSSd VDDd VSSd VSSd VSSd
+ VSSd VSSd SRegister_10_4/d SRegister_10_4/q out[6] out[4] out[10] out[7] out[5]
+ qw_NOLclk_0/PHI_2 out[8] VDDd SRegister_10_4/en VSSd qw_NOLclk_0/PHI_1 SRegister_10
Xasc_hysteresis_buffer_0 VSSd CLKd VDDd SCHMITT_0/IN asc_hysteresis_buffer
Xasc_hysteresis_buffer_1 VSSd ENd VDDd SRegister_10_4/en asc_hysteresis_buffer
Xasc_hysteresis_buffer_2 VSSd DATAd VDDd SRegister_10_4/d asc_hysteresis_buffer
XSCHMITT_0 VDDd VSSd SCHMITT_0/IN SCHMITT_0/OUT SCHMITT
XSRegister_10_0 out[31] out[32] out[33] out[39] VSSd VSSd VDDd VSSd VSSd VDDd VDDd
+ VSSd VSSd VSSd SRegister_10_3/q SRegister_10_2/d out[36] out[34] out[40] out[37]
+ out[35] qw_NOLclk_0/PHI_2 out[38] VDDd SRegister_10_4/en VSSd qw_NOLclk_0/PHI_1
+ SRegister_10
.ends

.subckt top_level_20250912_sc VDDd VSSd en clk data ref ext_pfd_div ext_pfd_ref ext_pfd_down
+ ext_pfd_up i_cp_100u up down lock filter_in filter_out ext_vco_in ext_vco_out out
+ div_in div_def div_out
Xtop_level_20250912_nosc_0 i_cp_100u div_def scan_chain_0/out[42] scan_chain_0/out[43]
+ scan_chain_0/out[44] scan_chain_0/out[45] scan_chain_0/out[46] scan_chain_0/out[47]
+ scan_chain_0/out[48] scan_chain_0/out[49] scan_chain_0/out[50] div_in scan_chain_0/out[41]
+ scan_chain_0/out[40] scan_chain_0/out[39] scan_chain_0/out[38] scan_chain_0/out[37]
+ scan_chain_0/out[36] scan_chain_0/out[35] scan_chain_0/out[34] scan_chain_0/out[33]
+ lock ref ext_pfd_div ext_pfd_ref ext_pfd_up ext_pfd_down scan_chain_0/out[1] scan_chain_0/out[2]
+ down scan_chain_0/out[6] scan_chain_0/out[5] scan_chain_0/out[4] scan_chain_0/out[3]
+ filter_in out filter_out scan_chain_0/out[32] scan_chain_0/out[31] scan_chain_0/out[26]
+ scan_chain_0/out[17] scan_chain_0/out[16] scan_chain_0/out[25] scan_chain_0/out[15]
+ scan_chain_0/out[24] scan_chain_0/out[14] scan_chain_0/out[13] scan_chain_0/out[12]
+ scan_chain_0/out[11] scan_chain_0/out[10] scan_chain_0/out[9] scan_chain_0/out[23]
+ scan_chain_0/out[22] scan_chain_0/out[21] scan_chain_0/out[20] scan_chain_0/out[19]
+ scan_chain_0/out[18] scan_chain_0/out[7] scan_chain_0/out[8] up ext_vco_out VDDd
+ VSSd ext_vco_in div_out top_level_20250912_nosc
Xscan_chain_0 VDDd en data clk scan_chain_0/out[1] scan_chain_0/out[2] scan_chain_0/out[3]
+ scan_chain_0/out[4] scan_chain_0/out[5] scan_chain_0/out[6] scan_chain_0/out[7]
+ scan_chain_0/out[8] scan_chain_0/out[9] scan_chain_0/out[10] scan_chain_0/out[20]
+ scan_chain_0/out[19] scan_chain_0/out[18] scan_chain_0/out[17] scan_chain_0/out[16]
+ scan_chain_0/out[15] scan_chain_0/out[14] scan_chain_0/out[13] scan_chain_0/out[12]
+ scan_chain_0/out[11] scan_chain_0/out[21] scan_chain_0/out[22] scan_chain_0/out[23]
+ scan_chain_0/out[24] scan_chain_0/out[25] scan_chain_0/out[26] scan_chain_0/out[27]
+ scan_chain_0/out[28] scan_chain_0/out[29] scan_chain_0/out[30] scan_chain_0/out[40]
+ scan_chain_0/out[39] scan_chain_0/out[38] scan_chain_0/out[37] scan_chain_0/out[36]
+ scan_chain_0/out[35] scan_chain_0/out[34] scan_chain_0/out[33] scan_chain_0/out[32]
+ scan_chain_0/out[31] scan_chain_0/out[41] scan_chain_0/out[42] scan_chain_0/out[43]
+ scan_chain_0/out[44] scan_chain_0/out[45] scan_chain_0/out[46] scan_chain_0/out[47]
+ scan_chain_0/out[48] scan_chain_0/out[49] scan_chain_0/out[50] VSSd scan_chain
.ends

