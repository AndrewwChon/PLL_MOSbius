* NGSPICE file created from xp_programmable_basic_pump.ext - technology: gf180mcuD

.subckt nfet$2 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$3 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_954_0# w_n180_n88# a_854_n136#
+ a_n92_0# a_446_n136# a_650_n136# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt pfet$1 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_954_0# w_n180_n88#
+ a_38_n60# a_n92_0# a_1058_n60# a_854_n60# a_342_0# a_138_0# a_650_n60#
X0 a_954_0# a_854_n60# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n60# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt pfet$7 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$6 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt inv1u05u VDD in VSS out w_2385_715# pfet$7_0/VSUBS
Xpfet$7_0 w_2385_715# VDD out in pfet$7
Xnfet$6_0 in VSS out pfet$7_0/VSUBS nfet$6
.ends

.subckt pfet$4 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.5u
.ends

.subckt pfet w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pass1u05u VDD clkp VSS clkn ins pfet_0/VSUBS w_3278_n1667# ind
Xpfet_0 w_3278_n1667# ind ins clkp pfet
Xnfet_0 clkn ind ins pfet_0/VSUBS nfet
.ends

.subckt pfet$2 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=4.55p ps=15.3u w=7u l=0.5u
.ends

.subckt nfet$5 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$1 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt nfet$2$1 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt xp_programmable_basic_pump VDD VSS up s1 s2 s3 s4 out iref down
Xnfet$2_2 VSS down VSS m1_592_n5360# down pfet$4_3/VSUBS nfet$2
Xnfet$2_15 m1_n774_n10170# pass1u05u_2/ins m1_n774_n10170# out pass1u05u_2/ins pfet$4_3/VSUBS
+ nfet$2
Xpfet$3_9 VDD VDD inv1u05u_0/out m3_1828_804# m3_1828_804# w_n10113_n2002# inv1u05u_0/out
+ VDD inv1u05u_0/out inv1u05u_0/out VDD m3_1828_804# inv1u05u_0/out inv1u05u_0/out
+ pfet$3
Xpfet$1_6 m3_851_5951# m3_851_5951# out pass1u05u_6/ins pass1u05u_6/ins out w_n10113_n2002#
+ pass1u05u_6/ins m3_851_5951# pass1u05u_6/ins pass1u05u_6/ins m3_851_5951# out pass1u05u_6/ins
+ pfet$1
Xinv1u05u_3 VDD s2 VSS inv1u05u_3/out w_4896_n9881# pfet$4_3/VSUBS inv1u05u
Xnfet$2_3 VSS down VSS m1_592_n5360# down pfet$4_3/VSUBS nfet$2
Xpfet$1_7 VDD VDD VDD VDD VDD VDD w_n10113_n2002# VDD VDD VDD VDD VDD VDD VDD pfet$1
Xinv1u05u_4 VDD s1 VSS inv1u05u_4/out w_4896_n9881# pfet$4_3/VSUBS inv1u05u
Xnfet$2_4 VSS down VSS m1_592_n5360# down pfet$4_3/VSUBS nfet$2
Xpfet$1_8 VDD VDD VDD VDD VDD VDD w_n10113_n2002# VDD VDD VDD VDD VDD VDD VDD pfet$1
Xnfet$2_5 VSS down VSS m1_592_n5360# down pfet$4_3/VSUBS nfet$2
Xpfet$1_9 m3_266_3959# m3_266_3959# pass1u05u_7/ind pass1u05u_7/ind pass1u05u_7/ind
+ pass1u05u_7/ind w_n10113_n2002# pass1u05u_7/ind m3_266_3959# pass1u05u_7/ind pass1u05u_7/ind
+ m3_266_3959# pass1u05u_7/ind pass1u05u_7/ind pfet$1
Xnfet$2_6 m1_592_n5360# pass1u05u_1/ins m1_592_n5360# out pass1u05u_1/ins pfet$4_3/VSUBS
+ nfet$2
Xnfet$2_7 m1_592_n5360# pass1u05u_1/ins m1_592_n5360# out pass1u05u_1/ins pfet$4_3/VSUBS
+ nfet$2
Xnfet$2_8 VSS down VSS m1_n774_n10170# down pfet$4_3/VSUBS nfet$2
Xnfet$2_9 VSS VDD VSS m3_n3965_n9526# VDD pfet$4_3/VSUBS nfet$2
Xpfet$4_0 w_4900_n7119# s3 pass1u05u_6/ins VDD pfet$4
Xpfet$4_1 w_4900_n7119# s2 pass1u05u_5/ins VDD pfet$4
Xpfet$4_2 w_4900_n7119# s1 pass1u05u_4/ins VDD pfet$4
Xpfet$4_3 w_4900_n7119# s4 pass1u05u_7/ins VDD pfet$4
Xpass1u05u_0 VDD inv1u05u_1/out VSS s4 pass1u05u_0/ins pfet$4_3/VSUBS w_4900_n7119#
+ iref pass1u05u
Xpfet$2_0 w_n10113_n2002# VDD VDD VDD pfet$2
Xnfet$5_0 inv1u05u_1/out pass1u05u_0/ins VSS pfet$4_3/VSUBS nfet$5
Xpass1u05u_1 VDD inv1u05u_2/out VSS s3 pass1u05u_1/ins pfet$4_3/VSUBS w_4900_n7119#
+ iref pass1u05u
Xpfet$2_1 w_n10113_n2002# VDD VDD VDD pfet$2
Xnfet$5_1 inv1u05u_2/out pass1u05u_1/ins VSS pfet$4_3/VSUBS nfet$5
Xpfet$2_10 w_n10113_n2002# VDD VDD VDD pfet$2
Xpfet$2_2 w_n10113_n2002# VDD VDD VDD pfet$2
Xpass1u05u_2 VDD inv1u05u_3/out VSS s2 pass1u05u_2/ins pfet$4_3/VSUBS w_4900_n7119#
+ iref pass1u05u
Xnfet$5_2 inv1u05u_3/out pass1u05u_2/ins VSS pfet$4_3/VSUBS nfet$5
Xpfet$2_11 w_n10113_n2002# VDD VDD VDD pfet$2
Xpfet$2_3 w_n10113_n2002# VDD VDD VDD pfet$2
Xpass1u05u_3 VDD inv1u05u_4/out VSS s1 pass1u05u_3/ins pfet$4_3/VSUBS w_4900_n7119#
+ iref pass1u05u
Xnfet$5_3 inv1u05u_4/out pass1u05u_3/ins VSS pfet$4_3/VSUBS nfet$5
Xpfet$2_4 w_n10113_n2002# VDD VDD VDD pfet$2
Xpass1u05u_4 VDD inv1u05u_4/out pass1u05u_7/VSS s1 pass1u05u_4/ins pfet$4_3/VSUBS
+ w_4900_n7119# pass1u05u_7/ind pass1u05u
Xpfet$2_5 w_n10113_n2002# VDD VDD VDD pfet$2
Xpass1u05u_5 VDD inv1u05u_3/out pass1u05u_7/VSS s2 pass1u05u_5/ins pfet$4_3/VSUBS
+ w_4900_n7119# pass1u05u_7/ind pass1u05u
Xpass1u05u_6 VDD inv1u05u_2/out pass1u05u_7/VSS s3 pass1u05u_6/ins pfet$4_3/VSUBS
+ w_4900_n7119# pass1u05u_7/ind pass1u05u
Xpfet$2_6 w_n10113_n2002# VDD VDD VDD pfet$2
Xnfet$1_0 VSS VSS VSS VSS VSS pfet$4_3/VSUBS nfet$1
Xpass1u05u_7 VDD inv1u05u_1/out pass1u05u_7/VSS s4 pass1u05u_7/ins pfet$4_3/VSUBS
+ w_4900_n7119# pass1u05u_7/ind pass1u05u
Xpfet$2_7 w_n10113_n2002# VDD VDD VDD pfet$2
Xnfet$1_1 VSS VSS VSS VSS VSS pfet$4_3/VSUBS nfet$1
Xpfet$2_8 w_n10113_n2002# VDD VDD VDD pfet$2
Xnfet$1_10 VSS VSS VSS VSS VSS pfet$4_3/VSUBS nfet$1
Xnfet$1_2 VSS VSS VSS VSS VSS pfet$4_3/VSUBS nfet$1
Xpfet$2_9 w_n10113_n2002# VDD VDD VDD pfet$2
Xnfet$1_11 pass1u05u_3/ins pass1u05u_3/ins m1_953_n7931# m1_953_n7931# out pfet$4_3/VSUBS
+ nfet$1
Xnfet$1_3 VSS VSS VSS VSS VSS pfet$4_3/VSUBS nfet$1
Xnfet$1_12 VSS VSS VSS VSS VSS pfet$4_3/VSUBS nfet$1
Xnfet$1_4 pass1u05u_0/ins pass1u05u_0/ins m1_n640_n5360# m1_n640_n5360# out pfet$4_3/VSUBS
+ nfet$1
Xnfet$1_13 down down VSS VSS m1_953_n7931# pfet$4_3/VSUBS nfet$1
Xnfet$1_5 pass1u05u_0/ins pass1u05u_0/ins m1_n640_n5360# m1_n640_n5360# out pfet$4_3/VSUBS
+ nfet$1
Xnfet$1_14 pass1u05u_0/ins pass1u05u_0/ins m1_n640_n5360# m1_n640_n5360# out pfet$4_3/VSUBS
+ nfet$1
Xnfet$1_6 pass1u05u_0/ins pass1u05u_0/ins m1_n640_n5360# m1_n640_n5360# out pfet$4_3/VSUBS
+ nfet$1
Xnfet$1_15 pass1u05u_0/ins pass1u05u_0/ins m1_n640_n5360# m1_n640_n5360# out pfet$4_3/VSUBS
+ nfet$1
Xpfet$3_20 m3_1828_804# m3_1828_804# pass1u05u_7/ins out out w_n10113_n2002# pass1u05u_7/ins
+ m3_1828_804# pass1u05u_7/ins pass1u05u_7/ins m3_1828_804# out pass1u05u_7/ins pass1u05u_7/ins
+ pfet$3
Xnfet$2$1_0 VSS VSS VSS VSS VSS pfet$4_3/VSUBS nfet$2$1
Xnfet$1_7 pass1u05u_0/ins pass1u05u_0/ins m1_n640_n5360# m1_n640_n5360# out pfet$4_3/VSUBS
+ nfet$1
Xpfet$3_21 m3_1828_804# m3_1828_804# pass1u05u_7/ins out out w_n10113_n2002# pass1u05u_7/ins
+ m3_1828_804# pass1u05u_7/ins pass1u05u_7/ins m3_1828_804# out pass1u05u_7/ins pass1u05u_7/ins
+ pfet$3
Xpfet$3_10 VDD VDD inv1u05u_0/out m3_851_5951# m3_851_5951# w_n10113_n2002# inv1u05u_0/out
+ VDD inv1u05u_0/out inv1u05u_0/out VDD m3_851_5951# inv1u05u_0/out inv1u05u_0/out
+ pfet$3
Xnfet$1_8 pass1u05u_0/ins pass1u05u_0/ins m1_n640_n5360# m1_n640_n5360# out pfet$4_3/VSUBS
+ nfet$1
Xnfet$2$1_1 down down VSS VSS m1_n640_n5360# pfet$4_3/VSUBS nfet$2$1
Xpfet$3_11 VDD VDD inv1u05u_0/out m3_266_4609# m3_266_4609# w_n10113_n2002# inv1u05u_0/out
+ VDD inv1u05u_0/out inv1u05u_0/out VDD m3_266_4609# inv1u05u_0/out inv1u05u_0/out
+ pfet$3
Xpfet$3_22 m3_1828_804# m3_1828_804# pass1u05u_7/ins out out w_n10113_n2002# pass1u05u_7/ins
+ m3_1828_804# pass1u05u_7/ins pass1u05u_7/ins m3_1828_804# out pass1u05u_7/ins pass1u05u_7/ins
+ pfet$3
Xnfet$1_9 pass1u05u_0/ins pass1u05u_0/ins m1_n640_n5360# m1_n640_n5360# out pfet$4_3/VSUBS
+ nfet$1
Xnfet$2$1_2 down down VSS VSS m1_n640_n5360# pfet$4_3/VSUBS nfet$2$1
Xpfet$3_12 VDD VDD inv1u05u_0/out m3_1476_2264# m3_1476_2264# w_n10113_n2002# inv1u05u_0/out
+ VDD inv1u05u_0/out inv1u05u_0/out VDD m3_1476_2264# inv1u05u_0/out inv1u05u_0/out
+ pfet$3
Xpfet$3_23 m3_266_4609# m3_266_4609# pass1u05u_4/ins out out w_n10113_n2002# pass1u05u_4/ins
+ m3_266_4609# pass1u05u_4/ins pass1u05u_4/ins m3_266_4609# out pass1u05u_4/ins pass1u05u_4/ins
+ pfet$3
Xpfet$3_0 VDD VDD inv1u05u_0/out m3_1828_804# m3_1828_804# w_n10113_n2002# inv1u05u_0/out
+ VDD inv1u05u_0/out inv1u05u_0/out VDD m3_1828_804# inv1u05u_0/out inv1u05u_0/out
+ pfet$3
Xnfet$2$1_10 down down VSS VSS m1_n640_n5360# pfet$4_3/VSUBS nfet$2$1
Xnfet$2$1_3 VSS VSS VSS VSS VSS pfet$4_3/VSUBS nfet$2$1
Xpfet$3_24 m3_1476_2264# m3_1476_2264# pass1u05u_5/ins out out w_n10113_n2002# pass1u05u_5/ins
+ m3_1476_2264# pass1u05u_5/ins pass1u05u_5/ins m3_1476_2264# out pass1u05u_5/ins
+ pass1u05u_5/ins pfet$3
Xpfet$3_13 VDD VDD inv1u05u_0/out m3_851_5951# m3_851_5951# w_n10113_n2002# inv1u05u_0/out
+ VDD inv1u05u_0/out inv1u05u_0/out VDD m3_851_5951# inv1u05u_0/out inv1u05u_0/out
+ pfet$3
Xpfet$3_1 VDD VDD inv1u05u_0/out m3_1828_804# m3_1828_804# w_n10113_n2002# inv1u05u_0/out
+ VDD inv1u05u_0/out inv1u05u_0/out VDD m3_1828_804# inv1u05u_0/out inv1u05u_0/out
+ pfet$3
Xnfet$2$1_11 down down VSS VSS m1_n640_n5360# pfet$4_3/VSUBS nfet$2$1
Xnfet$2$1_4 down down VSS VSS m1_n640_n5360# pfet$4_3/VSUBS nfet$2$1
Xpfet$3_25 m3_1476_2264# m3_1476_2264# pass1u05u_5/ins out out w_n10113_n2002# pass1u05u_5/ins
+ m3_1476_2264# pass1u05u_5/ins pass1u05u_5/ins m3_1476_2264# out pass1u05u_5/ins
+ pass1u05u_5/ins pfet$3
Xpfet$3_14 VDD VDD inv1u05u_0/out m3_1476_2264# m3_1476_2264# w_n10113_n2002# inv1u05u_0/out
+ VDD inv1u05u_0/out inv1u05u_0/out VDD m3_1476_2264# inv1u05u_0/out inv1u05u_0/out
+ pfet$3
Xpfet$3_2 VDD VDD inv1u05u_0/out m3_851_5951# m3_851_5951# w_n10113_n2002# inv1u05u_0/out
+ VDD inv1u05u_0/out inv1u05u_0/out VDD m3_851_5951# inv1u05u_0/out inv1u05u_0/out
+ pfet$3
Xnfet$2$1_12 VSS VSS VSS VSS VSS pfet$4_3/VSUBS nfet$2$1
Xnfet$2$1_5 down down VSS VSS m1_n640_n5360# pfet$4_3/VSUBS nfet$2$1
Xpfet$3_15 m3_1828_804# m3_1828_804# pass1u05u_7/ins out out w_n10113_n2002# pass1u05u_7/ins
+ m3_1828_804# pass1u05u_7/ins pass1u05u_7/ins m3_1828_804# out pass1u05u_7/ins pass1u05u_7/ins
+ pfet$3
Xpfet$3_3 VDD VDD inv1u05u_0/out m3_1828_804# m3_1828_804# w_n10113_n2002# inv1u05u_0/out
+ VDD inv1u05u_0/out inv1u05u_0/out VDD m3_1828_804# inv1u05u_0/out inv1u05u_0/out
+ pfet$3
Xnfet$2$1_13 VSS VSS VSS VSS VSS pfet$4_3/VSUBS nfet$2$1
Xpfet$1_0 VDD VDD VDD VDD VDD VDD w_n10113_n2002# VDD VDD VDD VDD VDD VDD VDD pfet$1
Xnfet$2$1_6 VSS VSS VSS VSS VSS pfet$4_3/VSUBS nfet$2$1
Xpfet$3_16 m3_1828_804# m3_1828_804# pass1u05u_7/ins out out w_n10113_n2002# pass1u05u_7/ins
+ m3_1828_804# pass1u05u_7/ins pass1u05u_7/ins m3_1828_804# out pass1u05u_7/ins pass1u05u_7/ins
+ pfet$3
Xnfet$2_10 m1_1576_n7920# iref m1_1576_n7920# pass1u05u_7/ind iref pfet$4_3/VSUBS
+ nfet$2
Xpfet$3_4 VDD VDD inv1u05u_0/out m3_1828_804# m3_1828_804# w_n10113_n2002# inv1u05u_0/out
+ VDD inv1u05u_0/out inv1u05u_0/out VDD m3_1828_804# inv1u05u_0/out inv1u05u_0/out
+ pfet$3
Xpfet$1_1 VDD VDD m3_266_3959# VSS VSS m3_266_3959# w_n10113_n2002# VSS VDD VSS VSS
+ VDD m3_266_3959# VSS pfet$1
Xnfet$2$1_7 VSS VSS VSS VSS VSS pfet$4_3/VSUBS nfet$2$1
Xpfet$3_17 m3_1828_804# m3_1828_804# pass1u05u_7/ins out out w_n10113_n2002# pass1u05u_7/ins
+ m3_1828_804# pass1u05u_7/ins pass1u05u_7/ins m3_1828_804# out pass1u05u_7/ins pass1u05u_7/ins
+ pfet$3
Xnfet$2_11 m1_n774_n10170# pass1u05u_2/ins m1_n774_n10170# out pass1u05u_2/ins pfet$4_3/VSUBS
+ nfet$2
Xpfet$3_5 VDD VDD inv1u05u_0/out m3_851_5951# m3_851_5951# w_n10113_n2002# inv1u05u_0/out
+ VDD inv1u05u_0/out inv1u05u_0/out VDD m3_851_5951# inv1u05u_0/out inv1u05u_0/out
+ pfet$3
Xpfet$1_2 VDD VDD VDD VDD VDD VDD w_n10113_n2002# VDD VDD VDD VDD VDD VDD VDD pfet$1
Xnfet$2$1_8 down down VSS VSS m1_n640_n5360# pfet$4_3/VSUBS nfet$2$1
Xpfet$3_18 m3_1828_804# m3_1828_804# pass1u05u_7/ins out out w_n10113_n2002# pass1u05u_7/ins
+ m3_1828_804# pass1u05u_7/ins pass1u05u_7/ins m3_1828_804# out pass1u05u_7/ins pass1u05u_7/ins
+ pfet$3
Xpfet$3_6 VDD VDD inv1u05u_0/out m3_1828_804# m3_1828_804# w_n10113_n2002# inv1u05u_0/out
+ VDD inv1u05u_0/out inv1u05u_0/out VDD m3_1828_804# inv1u05u_0/out inv1u05u_0/out
+ pfet$3
Xnfet$2_12 m3_n3965_n9526# iref m3_n3965_n9526# iref iref pfet$4_3/VSUBS nfet$2
Xpfet$1_3 m3_851_5951# m3_851_5951# out pass1u05u_6/ins pass1u05u_6/ins out w_n10113_n2002#
+ pass1u05u_6/ins m3_851_5951# pass1u05u_6/ins pass1u05u_6/ins m3_851_5951# out pass1u05u_6/ins
+ pfet$1
Xnfet$2$1_9 down down VSS VSS m1_n640_n5360# pfet$4_3/VSUBS nfet$2$1
Xinv1u05u_0 inv1u05u_0/VDD up VSS inv1u05u_0/out w_4896_n9881# pfet$4_3/VSUBS inv1u05u
Xpfet$3_19 m3_1828_804# m3_1828_804# pass1u05u_7/ins out out w_n10113_n2002# pass1u05u_7/ins
+ m3_1828_804# pass1u05u_7/ins pass1u05u_7/ins m3_1828_804# out pass1u05u_7/ins pass1u05u_7/ins
+ pfet$3
Xnfet$2_0 m1_592_n5360# pass1u05u_1/ins m1_592_n5360# out pass1u05u_1/ins pfet$4_3/VSUBS
+ nfet$2
Xpfet$3_7 VDD VDD inv1u05u_0/out m3_1828_804# m3_1828_804# w_n10113_n2002# inv1u05u_0/out
+ VDD inv1u05u_0/out inv1u05u_0/out VDD m3_1828_804# inv1u05u_0/out inv1u05u_0/out
+ pfet$3
Xnfet$2_13 VSS down VSS m1_n774_n10170# down pfet$4_3/VSUBS nfet$2
Xpfet$1_4 m3_851_5951# m3_851_5951# out pass1u05u_6/ins pass1u05u_6/ins out w_n10113_n2002#
+ pass1u05u_6/ins m3_851_5951# pass1u05u_6/ins pass1u05u_6/ins m3_851_5951# out pass1u05u_6/ins
+ pfet$1
Xinv1u05u_1 VDD s4 VSS inv1u05u_1/out w_4896_n9881# pfet$4_3/VSUBS inv1u05u
Xnfet$2_1 m1_592_n5360# pass1u05u_1/ins m1_592_n5360# out pass1u05u_1/ins pfet$4_3/VSUBS
+ nfet$2
Xpfet$3_8 VDD VDD inv1u05u_0/out m3_1828_804# m3_1828_804# w_n10113_n2002# inv1u05u_0/out
+ VDD inv1u05u_0/out inv1u05u_0/out VDD m3_1828_804# inv1u05u_0/out inv1u05u_0/out
+ pfet$3
Xnfet$2_14 VSS VDD VSS m1_1576_n7920# VDD pfet$4_3/VSUBS nfet$2
Xpfet$1_5 m3_851_5951# m3_851_5951# out pass1u05u_6/ins pass1u05u_6/ins out w_n10113_n2002#
+ pass1u05u_6/ins m3_851_5951# pass1u05u_6/ins pass1u05u_6/ins m3_851_5951# out pass1u05u_6/ins
+ pfet$1
Xinv1u05u_2 VDD s3 VSS inv1u05u_2/out w_4896_n9881# pfet$4_3/VSUBS inv1u05u
.ends

