* NGSPICE file created from top_level_20250919_wire.ext - technology: gf180mcuD

.subckt pfet$118 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$126 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$124 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$121 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$119 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$127 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$117 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$125 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$120 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$128 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_hysteresis_buffer$13 vss in vdd out
Xpfet$118_0 vdd vdd m1_884_42# m1_348_648# pfet$118
Xnfet$126_0 in vss m1_348_648# vss nfet$126
Xnfet$124_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$124
Xpfet$121_0 vdd vdd m1_884_42# m1_1156_42# pfet$121
Xpfet$119_0 vdd vdd m1_348_648# in pfet$119
Xnfet$127_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$127
Xpfet$117_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd
+ m1_884_42# m1_884_42# pfet$117
Xnfet$125_0 m1_348_648# vss m1_884_42# vss nfet$125
Xpfet$120_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$120
Xnfet$128_0 m1_1156_42# vss m1_884_42# vss nfet$128
.ends

.subckt pfet$60 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$64 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$61 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$65 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt xp_3_1_MUX$5 S0 S1 VDD VSS OUT_1 C_1 B_1 A_1
Xpfet$60_0 VDD A_1 m1_239_n318# m1_n432_458# pfet$60
Xpfet$60_1 VDD C_1 OUT_1 S1 pfet$60
Xpfet$60_2 VDD B_1 m1_239_n318# S0 pfet$60
Xpfet$60_3 VDD m1_239_n318# OUT_1 m1_n432_n1290# pfet$60
Xnfet$64_0 m1_n432_n1290# C_1 OUT_1 VSS nfet$64
Xnfet$64_1 m1_n432_458# B_1 m1_239_n318# VSS nfet$64
Xnfet$64_2 S1 m1_239_n318# OUT_1 VSS nfet$64
Xnfet$64_3 S0 A_1 m1_239_n318# VSS nfet$64
Xpfet$61_0 VDD VDD m1_n432_n1290# S1 pfet$61
Xpfet$61_1 VDD VDD m1_n432_458# S0 pfet$61
Xnfet$65_1 S0 VSS m1_n432_458# VSS nfet$65
Xnfet$65_0 S1 VSS m1_n432_n1290# VSS nfet$65
.ends

.subckt nfet$4 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$5 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$10 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$30 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$2 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$4 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$3 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$1 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$28 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$27 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$6 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$18 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$17 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$24 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$31 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$25 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$23 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$8 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$7 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$16 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$29 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$22 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$15 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$21 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$6 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$2 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$9 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$14 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$20 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$13 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$3 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$7 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$12 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$36 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$11 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$28 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$21 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$10 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$34 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$27 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$33 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$5 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$26 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$19 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$32 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$25 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$31 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$18 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$24 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$1 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$9 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$17 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$30 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$23 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$16 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$22 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$15 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$14 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$20 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$8 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$13 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$37 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$12 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$29 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$11 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$35 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$33 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$26 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$32 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$19 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_dual_psd_def_20250809$5 vdd vss pd1 pd2 pd3 pd4 pd5 pd6 pd7 pd8 pd9 fout
+ sd1 sd2 sd3 sd4 sd5 sd6 sd7 sd8 sd9 fin define
Xnfet$4_5 m1_649_17714# m1_649_17714# vss vss m1_6971_20470# vss nfet$4
Xnfet$5_69 m1_17851_17714# vss m1_17381_17714# vss nfet$5
Xnfet$5_58 m1_23007_17836# m1_23930_15778# m1_23109_16202# vss nfet$5
Xnfet$5_47 m1_22034_17714# vss m1_22624_17518# vss nfet$5
Xnfet$10_6 m1_n910_23922# vss m1_n290_24224# vss nfet$10
Xnfet$5_25 m1_2092_17836# m1_3372_16080# m1_2905_18030# vss nfet$5
Xnfet$5_14 m1_6116_17343# m1_8172_15778# m1_7555_16080# vss nfet$5
Xnfet$5_36 m1_n3064_17714# vss m1_n2474_17518# vss nfet$5
Xpfet$30_0 vdd m1_n6380_21786# m1_n6380_21786# m1_n5019_19550# m1_n5227_20152# m1_n5227_20152#
+ pfet$30
Xnfet$2_2 m1_n7513_20152# vss m1_4509_24346# vss nfet$2
Xnfet$2_59 m1_19644_25858# m1_20268_25662# m1_20005_23922# vss nfet$2
Xnfet$2_48 m1_18073_21786# vss m1_23827_25858# vss nfet$2
Xnfet$2_37 m1_11039_21786# vss m1_15461_25858# vss nfet$2
Xnfet$2_26 m1_7095_25858# m1_9180_25658# m1_9973_24542# vss nfet$2
Xnfet$2_15 m1_7232_25662# m1_7456_23922# m1_7720_24542# vss nfet$2
Xpfet$4_31 vdd m1_n2543_20130# m1_n2543_20130# m1_20407_19850# m1_19969_19550# m1_19969_19550#
+ pfet$4
Xpfet$4_20 vdd m1_n3822_21786# m1_n3822_21786# m1_14009_19550# m1_9015_17714# m1_9015_17714#
+ pfet$4
Xpfet$3_9 vdd m1_3871_22513# m1_3871_22513# m1_3471_22402# m1_4005_21786# m1_4005_21786#
+ pfet$3
Xpfet$1_6 vdd vdd m1_3536_25662# m1_3394_25858# pfet$1
Xnfet$28_7 m1_n3822_21786# m1_n3822_21786# m1_n4485_21904# m1_n4485_21904# m1_n3724_21430#
+ vss nfet$28
Xpfet$1_65 vdd vdd m1_18073_21786# m1_20126_25858# pfet$1
Xpfet$1_54 vdd vdd m1_24808_24224# m1_24188_23922# pfet$1
Xpfet$1_43 vdd vdd m1_12805_21786# pd5 pfet$1
Xpfet$1_32 vdd vdd m1_7720_24542# m1_8076_24224# pfet$1
Xpfet$1_21 vdd m1_7456_23922# m1_7720_24542# m1_7095_25858# pfet$1
Xpfet$1_10 vdd m1_8076_24224# m1_9180_25658# m1_7095_25858# pfet$1
Xpfet$27_6 vdd vdd m1_n4623_25487# fin pfet$27
Xpfet$1_98 vdd m1_30095_25658# m1_30888_24542# m1_28147_25662# pfet$1
Xpfet$1_87 vdd vdd m1_28147_25662# m1_28010_25858# pfet$1
Xpfet$1_76 vdd m1_20005_23922# m1_20269_24542# m1_19644_25858# pfet$1
Xnfet$6_9 m1_23356_21786# vss m1_23486_21590# vss nfet$6
Xpfet$18_2 vdd m1_32818_21586# m1_32818_21586# m1_33050_22344# m1_30256_22102# m1_30256_22102#
+ pfet$18
Xnfet$17_0 m1_31535_22102# m1_32818_21586# vss vss nfet$17
Xnfet$24_1 m1_n6433_17343# m1_n4377_15778# m1_n4994_16080# vss nfet$24
Xnfet$31_2 m1_n10933_25858# m1_n10309_25662# m1_n10572_23922# vss nfet$31
Xpfet$25_3 vdd vdd m1_n3651_26174# m1_n3541_23922# pfet$25
Xnfet$4_6 m1_n1133_19550# m1_n1133_19550# vss vss m1_n695_20470# vss nfet$4
Xnfet$10_7 m1_25107_21786# vss m1_32193_25858# vss nfet$10
Xnfet$5_59 m1_17851_17714# vss m1_20721_15778# vss nfet$5
Xnfet$5_48 m1_18824_17836# m1_20104_16080# m1_19637_18030# vss nfet$5
Xnfet$5_26 m1_5302_17714# vss m1_5892_17518# vss nfet$5
Xnfet$5_15 m1_5302_17714# vss m1_8172_15778# vss nfet$5
Xnfet$5_37 m1_n7513_20152# vss m1_n2605_16080# vss nfet$5
Xpfet$30_1 vdd vdd vdd m1_n5019_22344# m1_n4485_21904# m1_n4485_21904# pfet$30
Xpfet$23_0 vdd m1_n10309_25662# m1_n10572_23922# m1_n10796_25662# pfet$23
Xnfet$2_3 m1_488_21786# vss m1_2912_25858# vss nfet$2
Xnfet$2_49 m1_19781_25662# m1_20005_23922# m1_20269_24542# vss nfet$2
Xnfet$2_38 m1_n7513_20152# vss m1_12875_24346# vss nfet$2
Xnfet$2_27 m1_7577_25858# vss m1_7719_25662# vss nfet$2
Xnfet$2_16 m1_4005_21786# vss m1_7095_25858# vss nfet$2
Xpfet$4_32 vdd m1_n2543_20130# m1_n2543_20130# m1_21043_19550# m1_17381_17714# m1_17381_17714#
+ pfet$4
Xpfet$4_21 vdd vdd vdd m1_13373_19850# m1_15171_20152# m1_15171_20152# pfet$4
Xpfet$4_10 vdd vdd vdd m1_9856_19850# m1_11654_20152# m1_11654_20152# pfet$4
Xpfet$8_0 vdd vdd m1_n7401_15478# sd9 pfet$8
Xnfet$28_8 m1_9624_19404# m1_9624_19404# vss vss m1_n3724_21430# vss nfet$28
Xpfet$1_7 vdd vdd m1_7232_25662# m1_7095_25858# pfet$1
Xpfet$1_99 vdd vdd m1_26705_24542# m1_24309_25858# pfet$1
Xpfet$1_88 vdd vdd m1_28634_25662# m1_28492_25858# pfet$1
Xpfet$1_77 vdd vdd m1_20269_24542# m1_20625_24224# pfet$1
Xpfet$1_66 vdd vdd m1_15461_25858# m1_11039_21786# pfet$1
Xpfet$1_55 vdd m1_24451_25662# m1_24188_23922# m1_23964_25662# pfet$1
Xpfet$1_44 vdd m1_15943_25858# vdd m1_17546_25658# pfet$1
Xpfet$1_33 vdd vdd m1_7522_21786# m1_7577_25858# pfet$1
Xpfet$1_22 vdd vdd m1_3537_24542# m1_3893_24224# pfet$1
Xpfet$1_11 vdd vdd m1_7719_25662# m1_7577_25858# pfet$1
Xpfet$27_7 vdd vdd m1_n3541_23922# m1_n3184_24224# pfet$27
Xnfet$24_2 m1_n6274_17836# m1_n5351_15778# m1_n6172_16202# vss nfet$24
Xnfet$31_3 m1_n10796_25662# m1_n9952_24224# m1_n8848_25658# vss nfet$31
Xpfet$25_4 vdd m1_n10452_25858# vdd m1_n4362_24346# pfet$25
Xnfet$4_7 m1_n7383_17599# m1_n7383_17599# vss vss m1_n63_20470# vss nfet$4
Xnfet$10_8 m1_32193_25858# vss m1_32330_25662# vss nfet$10
Xnfet$5_49 m1_21564_17714# vss m1_18665_17343# vss nfet$5
Xpfet$7_10 vdd vdd m1_29239_20152# m1_26063_15478# pfet$7
Xnfet$5_27 m1_1119_17714# vss m1_3989_15778# vss nfet$5
Xnfet$5_16 m1_6275_17836# m1_7198_15778# m1_6377_16202# vss nfet$5
Xnfet$5_38 m1_n2250_17343# m1_n1989_16202# m1_n2474_17518# vss nfet$5
Xpfet$16_0 vdd vdd vdd m1_36073_22344# define define pfet$16
Xpfet$30_2 vdd m1_n5764_21786# m1_n5764_21786# m1_n5019_22344# m1_n5227_21418# m1_n5227_21418#
+ pfet$30
Xpfet$23_1 vdd m1_n9952_24224# m1_n8848_25658# m1_n10933_25858# pfet$23
Xnfet$2_4 m1_2912_25858# vss m1_3049_25662# vss nfet$2
Xnfet$29_10 vss vss m1_n4978_24224# vss nfet$29
Xnfet$2_39 pd4 vss m1_9288_21786# vss nfet$2
Xpfet$4_33 vdd m1_n3206_20274# m1_n3206_20274# m1_24560_19550# m1_21564_17714# m1_21564_17714#
+ pfet$4
Xpfet$4_22 vdd vdd vdd m1_14009_19550# m1_9331_15478# m1_9331_15478# pfet$4
Xnfet$2_28 m1_3394_25858# vss m1_4005_21786# vss nfet$2
Xnfet$2_17 m1_11639_23922# vss m1_12259_24224# vss nfet$2
Xpfet$4_11 vdd vdd vdd m1_10492_19550# m1_5148_15478# m1_5148_15478# pfet$4
Xpfet$8_1 vdd vdd m1_21880_15478# sd2 pfet$8
Xnfet$28_9 m1_n6380_21786# m1_n6380_21786# m1_n6839_21786# m1_n6839_21786# m1_n6282_21430#
+ vss nfet$28
Xpfet$1_8 vdd vdd m1_8076_24224# m1_7456_23922# pfet$1
Xpfet$1_89 vdd vdd m1_19839_21786# pd7 pfet$1
Xpfet$1_78 vdd m1_20269_24542# vdd m1_21241_24346# pfet$1
Xpfet$1_67 vdd m1_15822_23922# m1_16086_24542# m1_15461_25858# pfet$1
Xpfet$1_56 vdd m1_24808_24224# m1_25912_25658# m1_23827_25858# pfet$1
Xpfet$1_45 vdd vdd m1_16442_24224# m1_15822_23922# pfet$1
Xpfet$1_34 vdd m1_9180_25658# m1_9973_24542# m1_7232_25662# pfet$1
Xpfet$1_23 vdd m1_3537_24542# vdd m1_4509_24346# pfet$1
Xpfet$1_12 vdd m1_7577_25858# vdd m1_9180_25658# pfet$1
Xpfet$27_8 vdd vdd m1_n2567_23922# m1_n7320_25516# pfet$27
Xpfet$25_5 vdd vdd m1_n10308_24542# m1_n9952_24224# pfet$25
Xnfet$4_8 m1_27003_19550# m1_27003_19550# vss vss m1_27441_20470# vss nfet$4
Xnfet$24_3 m1_n6433_17343# m1_n6172_16202# m1_n6657_17518# vss nfet$24
Xnfet$31_4 m1_n4623_25487# m1_n2567_23922# m1_n3184_24224# vss nfet$31
Xnfet$10_9 m1_n7513_20152# vss m1_33790_24346# vss nfet$10
Xnfet$5_28 m1_1933_17343# vss m1_2092_17836# vss nfet$5
Xnfet$5_17 m1_649_17714# vss m1_n2250_17343# vss nfet$5
Xnfet$5_39 m1_n3064_17714# vss m1_n3534_17714# vss nfet$5
Xpfet$16_1 vdd m1_35837_22102# m1_35837_22102# m1_36073_22344# fout fout pfet$16
Xpfet$7_11 vdd vdd m1_18688_20152# m1_13514_15478# pfet$7
Xnfet$22_0 m1_4620_20152# m1_4620_20152# m1_2590_19404# m1_2590_19404# m1_3454_20470#
+ vss nfet$22
Xpfet$23_2 vdd m1_n4362_24346# m1_n4847_25662# m1_n4464_25980# pfet$23
Xnfet$2_5 m1_2912_25858# m1_3536_25662# m1_3273_23922# vss nfet$2
Xnfet$29_11 m1_n10452_25858# vss m1_n4847_25662# vss nfet$29
Xnfet$2_29 m1_15943_25858# vss m1_14556_21786# vss nfet$2
Xpfet$4_34 vdd m1_n3206_20274# m1_n3206_20274# m1_23924_19850# m1_23486_19550# m1_23486_19550#
+ pfet$4
Xpfet$4_23 vdd vdd vdd m1_16890_19850# m1_18688_20152# m1_18688_20152# pfet$4
Xnfet$2_18 m1_7095_25858# vss m1_7232_25662# vss nfet$2
Xpfet$4_12 vdd m1_6107_19404# m1_6107_19404# m1_6975_19550# m1_649_17714# m1_649_17714#
+ pfet$4
Xpfet$8_2 vdd vdd m1_26063_15478# sd1 pfet$8
Xpfet$1_9 vdd m1_7719_25662# m1_7456_23922# m1_7232_25662# pfet$1
Xpfet$1_79 vdd m1_17546_25658# m1_18339_24542# m1_15598_25662# pfet$1
Xpfet$1_68 vdd vdd m1_16086_24542# m1_16442_24224# pfet$1
Xpfet$1_57 vdd vdd m1_24451_25662# m1_24309_25858# pfet$1
Xpfet$1_46 vdd m1_16442_24224# m1_17546_25658# m1_15461_25858# pfet$1
Xpfet$1_35 vdd m1_7720_24542# vdd m1_8692_24346# pfet$1
Xpfet$1_24 vdd vdd m1_5790_24542# m1_3394_25858# pfet$1
Xpfet$1_13 vdd vdd m1_12259_24224# m1_11639_23922# pfet$1
Xpfet$27_9 vdd vdd m1_n4464_25980# m1_n4623_25487# pfet$27
Xnfet$4_9 m1_25747_17714# m1_25747_17714# vss vss m1_28073_20470# vss nfet$4
Xnfet$24_4 m1_27031_17343# m1_27292_16202# m1_26807_17518# vss nfet$24
Xnfet$31_5 m1_n4464_25980# m1_n3541_23922# m1_n4362_24346# vss nfet$31
Xpfet$25_6 vdd m1_n10308_24542# vdd m1_n9336_24346# pfet$25
Xnfet$5_29 m1_3372_16080# vss m1_3015_15778# vss nfet$5
Xnfet$5_18 m1_1119_17714# vss m1_649_17714# vss nfet$5
Xpfet$7_12 vdd vdd m1_15171_20152# m1_9331_15478# pfet$7
Xnfet$22_1 m1_1103_20152# m1_1103_20152# m1_n927_19404# m1_n927_19404# m1_n63_20470#
+ vss nfet$22
Xpfet$23_3 vdd m1_n3184_24224# m1_n3651_26174# m1_n4623_25487# pfet$23
Xnfet$15_0 m1_21456_22513# m1_21456_22513# m1_30256_19792# m1_30256_19792# m1_30492_20470#
+ vss nfet$15
Xnfet$2_6 m1_3049_25662# m1_3893_24224# m1_4997_25658# vss nfet$2
Xnfet$29_12 m1_n10452_25858# vss m1_n5571_25662# vss nfet$29
Xpfet$21_0 vdd vdd m1_n7513_20152# m1_35837_22102# pfet$21
Xnfet$2_19 m1_7456_23922# vss m1_8076_24224# vss nfet$2
Xpfet$4_35 vdd m1_n3822_21786# m1_n3822_21786# m1_13373_19850# m1_12935_19550# m1_12935_19550#
+ pfet$4
Xpfet$4_24 vdd m1_n1927_20274# m1_n1927_20274# m1_16890_19850# m1_16452_19550# m1_16452_19550#
+ pfet$4
Xpfet$4_13 vdd m1_n927_19404# m1_n927_19404# m1_n695_19850# m1_n1133_19550# m1_n1133_19550#
+ pfet$4
Xpfet$6_0 vdd vdd m1_n6274_17836# m1_n6433_17343# pfet$6
Xpfet$1_69 vdd vdd m1_12875_24346# m1_n7513_20152# pfet$1
Xpfet$1_58 vdd vdd m1_23964_25662# m1_23827_25858# pfet$1
Xpfet$1_47 vdd vdd m1_15943_25858# m1_17058_24346# pfet$1
Xpfet$1_36 vdd vdd m1_8692_24346# m1_n7513_20152# pfet$1
Xpfet$1_25 vdd vdd m1_4005_21786# m1_3394_25858# pfet$1
Xpfet$1_14 vdd vdd m1_11902_25662# m1_11760_25858# pfet$1
Xnfet$24_5 m1_27031_17343# m1_29087_15778# m1_28470_16080# vss nfet$24
Xnfet$31_6 m1_n4464_25980# m1_n3184_24224# m1_n3651_26174# vss nfet$31
Xpfet$25_7 vdd vdd m1_n10452_25858# m1_n4978_24224# pfet$25
Xpfet$2_90 vdd m1_19747_15778# m1_18926_16202# m1_18665_17343# pfet$2
Xnfet$9_0 m1_n3534_17714# vss m1_n6433_17343# vss nfet$9
Xpfet$7_13 vdd vdd m1_16452_19550# m1_13198_17714# pfet$7
Xnfet$5_19 m1_n7513_20152# vss m1_1578_16080# vss nfet$5
Xpfet$23_4 vdd m1_n2567_23922# m1_n3184_24224# m1_n4464_25980# pfet$23
Xnfet$15_1 m1_14422_22513# m1_14422_22513# m1_31535_19792# m1_31535_19792# m1_31771_20470#
+ vss nfet$15
Xnfet$2_7 m1_3049_25662# m1_3273_23922# m1_3537_24542# vss nfet$2
Xnfet$22_2 m1_n3218_15478# m1_n3218_15478# m1_2590_19404# m1_2590_19404# m1_2822_20470#
+ vss nfet$22
Xnfet$29_13 fin vss m1_n4623_25487# vss nfet$29
Xpfet$14_0 vdd vdd m1_n1263_21786# pd1 pfet$14
Xpfet$4_25 vdd vdd vdd m1_17526_19550# m1_13514_15478# m1_13514_15478# pfet$4
Xpfet$4_14 vdd m1_n927_19404# m1_n927_19404# m1_n59_19550# m1_n7383_17599# m1_n7383_17599#
+ pfet$4
Xpfet$6_1 vdd vdd m1_n4377_15778# m1_n7247_17714# pfet$6
Xpfet$1_59 vdd vdd m1_16322_21786# pd6 pfet$1
Xpfet$1_48 vdd m1_16085_25662# m1_15822_23922# m1_15598_25662# pfet$1
Xpfet$1_37 vdd vdd m1_9973_24542# m1_7577_25858# pfet$1
Xpfet$1_26 vdd m1_4997_25658# m1_5790_24542# m1_3049_25662# pfet$1
Xpfet$1_15 vdd m1_11902_25662# m1_11639_23922# m1_11415_25662# pfet$1
Xnfet$24_6 m1_27190_17836# m1_28113_15778# m1_27292_16202# vss nfet$24
Xnfet$31_7 m1_n4623_25487# m1_n4362_24346# m1_n4847_25662# vss nfet$31
Xpfet$2_91 vdd m1_24287_16080# m1_23820_18030# m1_22848_17343# pfet$2
Xpfet$2_80 vdd vdd m1_15564_15778# m1_15921_16080# pfet$2
Xpfet$7_14 vdd vdd m1_23486_19550# m1_21564_17714# pfet$7
Xnfet$9_1 m1_n7513_20152# vss m1_n6788_16080# vss nfet$9
Xnfet$15_2 m1_17939_22513# m1_17939_22513# vss vss m1_31771_20470# vss nfet$15
Xnfet$2_8 m1_3394_25858# vss m1_3536_25662# vss nfet$2
Xnfet$22_3 m1_8137_20152# m1_8137_20152# m1_6107_19404# m1_6107_19404# m1_6971_20470#
+ vss nfet$22
Xpfet$23_5 vdd m1_n10572_23922# m1_n10308_24542# m1_n10933_25858# pfet$23
Xpfet$14_1 vdd vdd m1_2254_21786# pd2 pfet$14
Xnfet$20_0 fout vss m1_35837_22102# vss nfet$20
Xpfet$4_26 vdd m1_n1927_20274# m1_n1927_20274# m1_17526_19550# m1_13198_17714# m1_13198_17714#
+ pfet$4
Xpfet$4_15 vdd vdd vdd m1_n59_19550# m1_n7401_15478# m1_n7401_15478# pfet$4
Xpfet$6_2 vdd vdd m1_n5351_15778# m1_n4994_16080# pfet$6
Xpfet$1_49 vdd m1_20126_25858# vdd m1_21729_25658# pfet$1
Xpfet$1_38 vdd vdd m1_16085_25662# m1_15943_25858# pfet$1
Xpfet$1_27 vdd vdd m1_11278_25858# m1_7522_21786# pfet$1
Xpfet$1_16 vdd vdd m1_5771_21786# pd3 pfet$1
Xnfet$24_7 m1_27190_17836# m1_28470_16080# m1_28003_18030# vss nfet$24
Xpfet$2_92 vdd m1_15454_18030# vdd m1_14127_16080# pfet$2
Xpfet$2_81 vdd vdd m1_13668_17714# m1_14127_16080# pfet$2
Xpfet$2_70 vdd vdd m1_18824_17836# m1_18665_17343# pfet$2
Xpfet$7_15 vdd vdd m1_22205_20152# m1_17697_15478# pfet$7
Xnfet$9_2 m1_n4994_16080# vss m1_n5351_15778# vss nfet$9
Xnfet$15_3 m1_24973_22513# m1_24973_22513# vss vss m1_30492_20470# vss nfet$15
Xnfet$22_4 m1_965_15478# m1_965_15478# m1_6107_19404# m1_6107_19404# m1_6339_20470#
+ vss nfet$22
Xpfet$23_6 vdd m1_n8848_25658# m1_n8055_24542# m1_n10796_25662# pfet$23
Xnfet$2_9 m1_3273_23922# vss m1_3893_24224# vss nfet$2
Xpfet$14_2 vdd vdd m1_26873_21786# pd9 pfet$14
Xnfet$20_1 define m1_35837_22102# vss vss nfet$20
Xnfet$13_0 m1_n290_24224# m1_n290_24224# m1_n646_24542# m1_n646_24542# m1_n192_24542#
+ vss nfet$13
Xpfet$4_27 vdd vdd vdd m1_20407_19850# m1_22205_20152# m1_22205_20152# pfet$4
Xpfet$4_16 vdd vdd vdd m1_28077_19550# m1_26063_15478# m1_26063_15478# pfet$4
Xnfet$3_10 m1_19839_21786# m1_19839_21786# m1_21456_22513# m1_21456_22513# m1_21060_21586#
+ vss nfet$3
Xpfet$6_3 vdd vdd m1_n6657_17518# m1_n7247_17714# pfet$6
Xpfet$1_39 vdd vdd m1_15598_25662# m1_15461_25858# pfet$1
Xpfet$1_28 vdd m1_11639_23922# m1_11903_24542# m1_11278_25858# pfet$1
Xpfet$1_17 vdd vdd m1_7577_25858# m1_8692_24346# pfet$1
Xpfet$4_0 vdd m1_2590_19404# m1_2590_19404# m1_3458_19550# m1_n3534_17714# m1_n3534_17714#
+ pfet$4
Xpfet$2_93 vdd m1_23820_18030# vdd m1_22493_16080# pfet$2
Xpfet$2_82 vdd m1_13668_17714# vdd m1_14743_16202# pfet$2
Xpfet$2_71 vdd vdd m1_19747_15778# m1_20104_16080# pfet$2
Xpfet$2_60 vdd vdd m1_n194_15778# m1_n3064_17714# pfet$2
Xnfet$9_3 m1_n6433_17343# vss m1_n6274_17836# vss nfet$9
Xpfet$7_16 vdd vdd m1_19969_19550# m1_17381_17714# pfet$7
Xnfet$15_4 m1_32818_20470# m1_32818_20470# vss vss m1_34329_20470# vss nfet$15
Xnfet$22_5 m1_5148_15478# m1_5148_15478# m1_9624_19404# m1_9624_19404# m1_9856_20470#
+ vss nfet$22
Xpfet$23_7 vdd m1_n3541_23922# m1_n4362_24346# m1_n4623_25487# pfet$23
Xnfet$7_0 m1_n3534_17714# vss m1_2384_19550# vss nfet$7
Xnfet$6_10 m1_21590_21786# vss m1_22222_21786# vss nfet$6
Xnfet$13_1 m1_814_25658# m1_814_25658# vss vss m1_1273_25502# vss nfet$13
Xpfet$4_28 vdd vdd vdd m1_21043_19550# m1_17697_15478# m1_17697_15478# pfet$4
Xpfet$4_17 vdd m1_n3822_20130# m1_n3822_20130# m1_28077_19550# m1_25747_17714# m1_25747_17714#
+ pfet$4
Xpfet$12_0 vdd m1_31535_19792# vdd m1_17939_22513# pfet$12
Xnfet$3_11 m1_19969_21590# m1_19969_21590# m1_21456_22513# m1_21456_22513# m1_20428_21586#
+ vss nfet$3
Xpfet$6_4 vdd vdd m1_n6433_17343# m1_n3534_17714# pfet$6
Xpfet$1_29 vdd vdd m1_11903_24542# m1_12259_24224# pfet$1
Xpfet$1_18 vdd vdd m1_11415_25662# m1_11278_25858# pfet$1
Xpfet$4_1 vdd vdd vdd m1_2822_19850# m1_4620_20152# m1_4620_20152# pfet$4
Xnfet$9_10 m1_26217_17714# vss m1_29087_15778# vss nfet$9
Xpfet$2_94 vdd vdd m1_22624_17518# m1_22034_17714# pfet$2
Xpfet$2_83 vdd m1_16538_15778# m1_15921_16080# m1_14641_17836# pfet$2
Xpfet$2_72 vdd m1_20721_15778# m1_20104_16080# m1_18824_17836# pfet$2
Xpfet$2_61 vdd m1_n811_16080# m1_n1278_18030# m1_n2250_17343# pfet$2
Xpfet$2_50 vdd m1_n1168_15778# m1_n1989_16202# m1_n2250_17343# pfet$2
Xnfet$9_4 m1_n7247_17714# vss m1_n4377_15778# vss nfet$9
Xnfet$36_0 m1_n4485_20152# m1_n6380_21786# vss vss nfet$36
Xpfet$7_17 vdd vdd m1_25722_20152# m1_21880_15478# pfet$7
Xnfet$22_6 m1_11654_20152# m1_11654_20152# m1_9624_19404# m1_9624_19404# m1_10488_20470#
+ vss nfet$22
Xnfet$15_5 m1_32818_21586# m1_32818_21586# m1_34093_19792# m1_34093_19792# m1_34329_20470#
+ vss nfet$15
Xnfet$7_1 m1_n3218_15478# vss m1_4620_20152# vss nfet$7
Xnfet$6_11 m1_18073_21786# vss m1_18705_21786# vss nfet$6
Xnfet$13_2 m1_326_24346# m1_326_24346# m1_n789_25858# m1_n789_25858# m1_1273_25502#
+ vss nfet$13
Xpfet$4_29 vdd vdd vdd m1_23924_19850# m1_25722_20152# m1_25722_20152# pfet$4
Xpfet$4_18 vdd vdd vdd m1_27441_19850# m1_29239_20152# m1_29239_20152# pfet$4
Xpfet$12_1 vdd vdd m1_30256_19792# m1_21456_22513# pfet$12
Xnfet$3_12 m1_16322_21786# m1_16322_21786# m1_17939_22513# m1_17939_22513# m1_17543_21586#
+ vss nfet$3
Xpfet$6_5 vdd vdd m1_n6788_16080# m1_n7513_20152# pfet$6
Xpfet$1_19 vdd vdd m1_7095_25858# m1_4005_21786# pfet$1
Xpfet$4_2 vdd m1_2590_19404# m1_2590_19404# m1_2822_19850# m1_2384_19550# m1_2384_19550#
+ pfet$4
Xnfet$9_11 m1_27031_17343# vss m1_27190_17836# vss nfet$9
Xpfet$2_95 vdd vdd m1_21564_17714# m1_22034_17714# pfet$2
Xpfet$2_84 vdd vdd m1_17381_17714# m1_17851_17714# pfet$2
Xpfet$2_73 vdd vdd m1_16538_15778# m1_13668_17714# pfet$2
Xpfet$2_62 vdd vdd m1_23007_17836# m1_22848_17343# pfet$2
Xpfet$2_40 vdd m1_10560_16202# m1_10075_17518# m1_10458_17836# pfet$2
Xpfet$2_51 vdd vdd m1_n1168_15778# m1_n811_16080# pfet$2
Xnfet$9_5 m1_n7247_17714# vss m1_n6657_17518# vss nfet$9
Xnfet$36_1 m1_n5227_20152# vss m1_n6380_21786# vss nfet$36
Xnfet$29_0 m1_n8625_26174# vss m1_n8055_24542# vss nfet$29
Xnfet$15_6 m1_354_22513# m1_354_22513# m1_31535_22102# m1_31535_22102# m1_31771_21430#
+ vss nfet$15
Xnfet$22_7 m1_n7401_15478# m1_n7401_15478# m1_n927_19404# m1_n927_19404# m1_n695_20470#
+ vss nfet$22
Xnfet$7_2 m1_n7401_15478# vss m1_1103_20152# vss nfet$7
Xnfet$6_12 m1_14556_21786# vss m1_15188_21786# vss nfet$6
Xnfet$13_3 m1_326_24346# m1_326_24346# vss vss m1_n192_24542# vss nfet$13
Xpfet$4_19 vdd m1_n3822_20130# m1_n3822_20130# m1_27441_19850# m1_27003_19550# m1_27003_19550#
+ pfet$4
Xpfet$12_2 vdd m1_30256_19792# vdd m1_24973_22513# pfet$12
Xnfet$11_0 m1_n1134_25662# m1_n910_23922# m1_n646_24542# vss nfet$11
Xnfet$3_13 m1_16452_21590# m1_16452_21590# m1_17939_22513# m1_17939_22513# m1_16911_21586#
+ vss nfet$3
Xpfet$6_6 vdd vdd m1_n7383_17599# m1_n7247_17714# pfet$6
Xpfet$4_3 vdd vdd vdd m1_3458_19550# m1_n3218_15478# m1_n3218_15478# pfet$4
Xpfet$2_96 vdd vdd m1_18665_17343# m1_21564_17714# pfet$2
Xpfet$2_85 vdd m1_18926_16202# m1_18441_17518# m1_18824_17836# pfet$2
Xpfet$2_74 vdd vdd m1_14641_17836# m1_14482_17343# pfet$2
Xpfet$2_63 vdd m1_23930_15778# m1_23109_16202# m1_22848_17343# pfet$2
Xnfet$9_12 m1_28470_16080# vss m1_28113_15778# vss nfet$9
Xpfet$2_30 vdd vdd m1_1933_17343# m1_4832_17714# pfet$2
Xpfet$2_41 vdd vdd m1_10075_17518# m1_9485_17714# pfet$2
Xpfet$2_52 vdd m1_n3064_17714# vdd m1_n1989_16202# pfet$2
Xnfet$29_1 m1_n8625_26174# vss m1_n7082_23622# vss nfet$29
Xpfet$2_0 vdd vdd m1_12355_15778# m1_9485_17714# pfet$2
Xnfet$9_6 m1_n7247_17714# vss m1_n7383_17599# vss nfet$9
Xnfet$15_7 m1_3871_22513# m1_3871_22513# vss vss m1_31771_21430# vss nfet$15
Xnfet$22_8 m1_26063_15478# m1_26063_15478# m1_n3822_20130# m1_n3822_20130# m1_27441_20470#
+ vss nfet$22
Xnfet$10_10 m1_32675_25947# vss m1_35071_24542# vss nfet$10
Xnfet$7_3 m1_649_17714# vss m1_5901_19550# vss nfet$7
Xpfet$28_0 vdd vdd m1_n7186_25858# m1_n10452_25858# pfet$28
Xnfet$6_13 m1_16322_21786# vss m1_16452_21590# vss nfet$6
Xnfet$13_4 m1_33174_24224# m1_33174_24224# m1_32818_24542# m1_32818_24542# m1_33272_24542#
+ vss nfet$13
Xnfet$21_20 m1_22493_16080# m1_22493_16080# m1_22034_17714# m1_22034_17714# m1_22591_16398#
+ vss nfet$21
Xnfet$5_0 m1_9485_17714# vss m1_9015_17714# vss nfet$5
Xpfet$12_3 vdd vdd m1_34843_21786# m1_34093_19792# pfet$12
Xnfet$11_1 m1_n1271_25858# m1_n647_25662# m1_n910_23922# vss nfet$11
Xnfet$3_14 m1_12805_21786# m1_12805_21786# m1_14422_22513# m1_14422_22513# m1_14026_21586#
+ vss nfet$3
Xpfet$6_7 vdd vdd m1_27190_17836# m1_27031_17343# pfet$6
Xpfet$10_0 vdd vdd m1_n646_24542# m1_n290_24224# pfet$10
Xpfet$4_4 vdd m1_6107_19404# m1_6107_19404# m1_6339_19850# m1_5901_19550# m1_5901_19550#
+ pfet$4
Xnfet$9_13 m1_26217_17714# vss m1_25747_17714# vss nfet$9
Xpfet$2_97 vdd vdd m1_22493_16080# m1_n7513_20152# pfet$2
Xpfet$2_86 vdd m1_19637_18030# vdd m1_18310_16080# pfet$2
Xpfet$2_75 vdd vdd m1_17697_15478# sd3 pfet$2
Xpfet$2_64 vdd vdd m1_23930_15778# m1_24287_16080# pfet$2
Xpfet$2_20 vdd vdd m1_1119_17714# m1_1578_16080# pfet$2
Xpfet$2_31 vdd m1_3372_16080# m1_2905_18030# m1_1933_17343# pfet$2
Xpfet$2_42 vdd m1_11271_18030# vdd m1_9944_16080# pfet$2
Xpfet$2_53 vdd vdd m1_n3218_15478# sd8 pfet$2
Xnfet$29_2 vss vss m1_n9336_24346# vss nfet$29
Xnfet$9_7 m1_26217_17714# vss m1_26807_17518# vss nfet$9
Xpfet$2_1 vdd vdd m1_11381_15778# m1_11738_16080# pfet$2
Xnfet$22_9 m1_29239_20152# m1_29239_20152# m1_n3822_20130# m1_n3822_20130# m1_28073_20470#
+ vss nfet$22
Xnfet$10_11 m1_32554_23922# vss m1_33174_24224# vss nfet$10
Xnfet$34_0 m1_n4485_21904# m1_n5764_21786# vss vss nfet$34
Xpfet$28_1 vdd m1_n7186_25858# vdd m1_n6111_25858# pfet$28
Xnfet$6_14 m1_19839_21786# vss m1_19969_21590# vss nfet$6
Xnfet$7_4 m1_4832_17714# vss m1_9418_19550# vss nfet$7
Xnfet$13_5 m1_33790_24346# m1_33790_24346# vss vss m1_33272_24542# vss nfet$13
Xnfet$21_21 m1_14127_16080# m1_14127_16080# vss vss m1_15690_17358# vss nfet$21
Xnfet$21_10 m1_1578_16080# m1_1578_16080# m1_1119_17714# m1_1119_17714# m1_1676_16398#
+ vss nfet$21
Xnfet$5_1 m1_9015_17714# vss m1_6116_17343# vss nfet$5
Xpfet$12_4 vdd m1_34093_19792# vdd m1_32818_20470# pfet$12
Xnfet$11_2 m1_n1271_25858# m1_814_25658# m1_1607_24542# vss nfet$11
Xnfet$3_15 m1_26873_21786# m1_26873_21786# m1_28490_22513# m1_28490_22513# m1_28094_21586#
+ vss nfet$3
Xpfet$6_8 vdd vdd m1_28113_15778# m1_28470_16080# pfet$6
Xpfet$10_1 vdd m1_n789_25858# vdd m1_814_25658# pfet$10
Xpfet$4_5 vdd vdd vdd m1_n695_19850# m1_1103_20152# m1_1103_20152# pfet$4
Xpfet$2_98 vdd m1_20104_16080# m1_19637_18030# m1_18665_17343# pfet$2
Xpfet$2_87 vdd vdd m1_18310_16080# m1_n7513_20152# pfet$2
Xpfet$2_76 vdd m1_17851_17714# vdd m1_18926_16202# pfet$2
Xpfet$2_65 vdd m1_24904_15778# m1_24287_16080# m1_23007_17836# pfet$2
Xpfet$2_21 vdd vdd m1_965_15478# sd7 pfet$2
Xpfet$2_10 vdd m1_8172_15778# m1_7555_16080# m1_6275_17836# pfet$2
Xpfet$2_32 vdd vdd m1_2905_18030# m1_3015_15778# pfet$2
Xpfet$2_43 vdd vdd m1_11271_18030# m1_11381_15778# pfet$2
Xpfet$2_54 vdd vdd m1_n1278_18030# m1_n1168_15778# pfet$2
Xnfet$29_3 fin vss m1_n10933_25858# vss nfet$29
Xnfet$9_8 m1_n7513_20152# vss m1_26676_16080# vss nfet$9
Xpfet$2_2 vdd m1_12355_15778# m1_11738_16080# m1_10458_17836# pfet$2
Xnfet$10_12 m1_32675_25947# vss m1_28624_21786# vss nfet$10
Xnfet$34_1 m1_n5227_21418# vss m1_n5764_21786# vss nfet$34
Xnfet$27_0 m1_n7082_23622# m1_n6856_24542# vss vss nfet$27
Xnfet$7_5 m1_965_15478# vss m1_8137_20152# vss nfet$7
Xnfet$13_6 m1_33790_24346# m1_33790_24346# m1_32675_25947# m1_32675_25947# m1_34737_25502#
+ vss nfet$13
Xnfet$6_15 m1_28624_21786# vss m1_29256_21786# vss nfet$6
Xnfet$21_22 m1_15564_15778# m1_15564_15778# m1_15454_18030# m1_15454_18030# m1_15690_17358#
+ vss nfet$21
Xnfet$5_2 m1_6275_17836# m1_7555_16080# m1_7088_18030# vss nfet$5
Xnfet$21_11 m1_6377_16202# m1_6377_16202# vss vss m1_5859_16398# vss nfet$21
Xpfet$33_0 vdd vdd m1_n8145_21908# m1_n6839_20152# pfet$33
Xpfet$12_5 vdd vdd m1_34093_19792# m1_32818_21586# pfet$12
Xnfet$11_3 m1_n1134_25662# m1_n290_24224# m1_814_25658# vss nfet$11
Xnfet$3_16 m1_27003_21590# m1_27003_21590# m1_28490_22513# m1_28490_22513# m1_27462_21586#
+ vss nfet$3
Xpfet$5_10 vdd vdd m1_23486_21590# m1_23356_21786# pfet$5
Xpfet$6_9 vdd vdd m1_29087_15778# m1_26217_17714# pfet$6
Xpfet$10_2 vdd vdd m1_n789_25858# m1_326_24346# pfet$10
Xpfet$4_6 vdd vdd vdd m1_6339_19850# m1_8137_20152# m1_8137_20152# pfet$4
Xpfet$2_22 vdd vdd m1_3015_15778# m1_3372_16080# pfet$2
Xpfet$2_11 vdd vdd m1_9485_17714# m1_9944_16080# pfet$2
Xpfet$2_33 vdd vdd m1_5892_17518# m1_5302_17714# pfet$2
Xpfet$2_99 vdd m1_23109_16202# m1_22624_17518# m1_23007_17836# pfet$2
Xpfet$2_88 vdd vdd m1_18441_17518# m1_17851_17714# pfet$2
Xpfet$2_77 vdd vdd m1_17851_17714# m1_18310_16080# pfet$2
Xpfet$2_66 vdd vdd m1_24904_15778# m1_22034_17714# pfet$2
Xnfet$9_9 m1_n10452_25858# vss m1_27031_17343# vss nfet$9
Xpfet$2_3 vdd m1_11381_15778# m1_10560_16202# m1_10299_17343# pfet$2
Xpfet$2_44 vdd vdd m1_649_17714# m1_1119_17714# pfet$2
Xpfet$2_55 vdd vdd m1_n2474_17518# m1_n3064_17714# pfet$2
Xnfet$29_4 m1_n10572_23922# vss m1_n9952_24224# vss nfet$29
Xnfet$34_2 m1_n6839_21786# vss m1_n6973_21481# vss nfet$34
Xnfet$27_1 m1_n8283_19850# vss m1_n6856_24542# vss nfet$27
Xnfet$10_13 m1_32675_25947# vss m1_32817_25662# vss nfet$10
Xnfet$7_6 m1_9015_17714# vss m1_12935_19550# vss nfet$7
Xpfet$2_110 vdd vdd m1_10458_17836# m1_10299_17343# pfet$2
Xnfet$13_7 m1_34278_25658# m1_34278_25658# vss vss m1_34737_25502# vss nfet$13
Xnfet$6_16 m1_26873_21786# vss m1_27003_21590# vss nfet$6
Xnfet$21_23 m1_18926_16202# m1_18926_16202# vss vss m1_18408_16398# vss nfet$21
Xnfet$21_12 m1_n1168_15778# m1_n1168_15778# m1_n1278_18030# m1_n1278_18030# m1_n1042_17358#
+ vss nfet$21
Xpfet$26_0 vdd vdd m1_n4485_20152# m1_n3822_20130# pfet$26
Xnfet$5_3 m1_n7513_20152# vss m1_9944_16080# vss nfet$5
Xnfet$11_4 m1_32193_25858# m1_34278_25658# m1_35071_24542# vss nfet$11
Xpfet$12_6 vdd vdd m1_31535_19792# m1_14422_22513# pfet$12
Xnfet$3_17 m1_12935_21590# m1_12935_21590# m1_14422_22513# m1_14422_22513# m1_13394_21586#
+ vss nfet$3
Xnfet$3_0 m1_n1133_21590# m1_n1133_21590# m1_354_22513# m1_354_22513# m1_n674_21586#
+ vss nfet$3
Xpfet$5_11 vdd vdd m1_18705_21786# m1_18073_21786# pfet$5
Xpfet$10_3 vdd m1_n646_24542# vdd m1_326_24346# pfet$10
Xpfet$4_7 vdd vdd vdd m1_6975_19550# m1_965_15478# m1_965_15478# pfet$4
Xpfet$2_89 vdd vdd m1_22848_17343# m1_25747_17714# pfet$2
Xpfet$2_78 vdd vdd m1_13514_15478# sd4 pfet$2
Xpfet$2_67 vdd m1_22034_17714# vdd m1_23109_16202# pfet$2
Xpfet$2_12 vdd m1_3989_15778# m1_3372_16080# m1_2092_17836# pfet$2
Xpfet$2_4 vdd m1_9485_17714# vdd m1_10560_16202# pfet$2
Xpfet$2_23 vdd m1_5302_17714# vdd m1_6377_16202# pfet$2
Xpfet$2_34 vdd vdd m1_5761_16080# m1_n7513_20152# pfet$2
Xpfet$2_45 vdd vdd m1_9944_16080# m1_n7513_20152# pfet$2
Xpfet$2_56 vdd m1_n1278_18030# vdd m1_n2605_16080# pfet$2
Xnfet$29_5 m1_n10933_25858# vss m1_n10796_25662# vss nfet$29
Xnfet$7_7 m1_5148_15478# vss m1_11654_20152# vss nfet$7
Xnfet$6_17 m1_25107_21786# vss m1_25739_21786# vss nfet$6
Xpfet$2_100 vdd vdd m1_23820_18030# m1_23930_15778# pfet$2
Xnfet$21_24 m1_18310_16080# m1_18310_16080# m1_17851_17714# m1_17851_17714# m1_18408_16398#
+ vss nfet$21
Xnfet$21_13 m1_n2605_16080# m1_n2605_16080# vss vss m1_n1042_17358# vss nfet$21
Xpfet$19_0 vdd vdd m1_n7247_17714# m1_n6788_16080# pfet$19
Xpfet$26_1 vdd m1_n4485_21904# vdd m1_9624_19404# pfet$26
Xnfet$32_0 m1_n7186_25858# vss m1_n7320_25516# vss nfet$32
Xnfet$5_4 m1_10299_17343# m1_10560_16202# m1_10075_17518# vss nfet$5
Xpfet$12_7 vdd vdd m1_31535_22102# m1_354_22513# pfet$12
Xnfet$11_5 m1_32330_25662# m1_33174_24224# m1_34278_25658# vss nfet$11
Xnfet$3_1 m1_n1263_21786# m1_n1263_21786# m1_354_22513# m1_354_22513# m1_n42_21586#
+ vss nfet$3
Xpfet$5_12 vdd vdd m1_16452_21590# m1_16322_21786# pfet$5
Xpfet$10_4 vdd vdd m1_32675_25947# m1_33790_24346# pfet$10
Xpfet$4_8 vdd m1_9624_19404# m1_9624_19404# m1_10492_19550# m1_4832_17714# m1_4832_17714#
+ pfet$4
Xpfet$2_79 vdd m1_15564_15778# m1_14743_16202# m1_14482_17343# pfet$2
Xpfet$2_68 vdd vdd m1_22034_17714# m1_22493_16080# pfet$2
Xpfet$2_13 vdd vdd m1_5148_15478# sd6 pfet$2
Xpfet$2_24 vdd m1_6377_16202# m1_5892_17518# m1_6275_17836# pfet$2
Xpfet$2_35 vdd vdd m1_9015_17714# m1_9485_17714# pfet$2
Xpfet$2_46 vdd vdd m1_n2250_17343# m1_649_17714# pfet$2
Xpfet$2_57 vdd m1_n1989_16202# m1_n2474_17518# m1_n2091_17836# pfet$2
Xnfet$29_6 m1_n10452_25858# vss m1_n10309_25662# vss nfet$29
Xpfet$2_5 vdd m1_7198_15778# m1_6377_16202# m1_6116_17343# pfet$2
Xnfet$7_8 m1_n7383_17599# vss m1_n1133_19550# vss nfet$7
Xpfet$2_101 vdd vdd m1_19637_18030# m1_19747_15778# pfet$2
Xnfet$25_0 m1_n5351_15778# m1_n5351_15778# m1_n5461_18030# m1_n5461_18030# m1_n5225_17358#
+ vss nfet$25
Xpfet$19_1 vdd m1_n7247_17714# vdd m1_n6172_16202# pfet$19
Xpfet$26_2 vdd m1_n5227_21418# vdd m1_2590_19404# pfet$26
Xnfet$32_1 m1_n6856_24542# vss m1_n6111_25858# vss nfet$32
Xnfet$21_25 m1_14743_16202# m1_14743_16202# vss vss m1_14225_16398# vss nfet$21
Xnfet$5_5 m1_10458_17836# m1_11738_16080# m1_11271_18030# vss nfet$5
Xnfet$21_14 m1_n2605_16080# m1_n2605_16080# m1_n3064_17714# m1_n3064_17714# m1_n2507_16398#
+ vss nfet$21
Xnfet$11_6 m1_32193_25858# m1_32817_25662# m1_32554_23922# vss nfet$11
Xpfet$31_0 vdd vdd m1_n5227_20152# m1_n2543_20130# pfet$31
Xpfet$5_13 vdd vdd m1_15188_21786# m1_14556_21786# pfet$5
Xnfet$3_2 m1_9288_21786# m1_9288_21786# m1_9645_21447# m1_9645_21447# m1_10509_21586#
+ vss nfet$3
Xpfet$10_5 vdd m1_32675_25947# vdd m1_34278_25658# pfet$10
Xpfet$4_9 vdd m1_9624_19404# m1_9624_19404# m1_9856_19850# m1_9418_19550# m1_9418_19550#
+ pfet$4
Xpfet$2_69 vdd vdd m1_20721_15778# m1_17851_17714# pfet$2
Xpfet$2_14 vdd vdd m1_2092_17836# m1_1933_17343# pfet$2
Xpfet$2_25 vdd vdd m1_1709_17518# m1_1119_17714# pfet$2
Xpfet$2_36 vdd vdd m1_6116_17343# m1_9015_17714# pfet$2
Xpfet$2_47 vdd m1_11738_16080# m1_11271_18030# m1_10299_17343# pfet$2
Xpfet$2_58 vdd vdd m1_n3534_17714# m1_n3064_17714# pfet$2
Xnfet$29_7 m1_n7320_25516# vss m1_n2567_23922# vss nfet$29
Xpfet$2_6 vdd vdd m1_7198_15778# m1_7555_16080# pfet$2
Xnfet$7_9 m1_25747_17714# vss m1_27003_19550# vss nfet$7
Xpfet$2_102 vdd vdd m1_13198_17714# m1_13668_17714# pfet$2
Xpfet$19_2 vdd vdd m1_n5461_18030# m1_n5351_15778# pfet$19
Xpfet$26_3 vdd vdd m1_n5227_21418# m1_6107_19404# pfet$26
Xnfet$21_26 m1_14127_16080# m1_14127_16080# m1_13668_17714# m1_13668_17714# m1_14225_16398#
+ vss nfet$21
Xnfet$18_0 m1_34093_19792# vss m1_34843_21786# vss nfet$18
Xnfet$5_6 m1_6116_17343# vss m1_6275_17836# vss nfet$5
Xnfet$25_1 m1_n6788_16080# m1_n6788_16080# vss vss m1_n5225_17358# vss nfet$25
Xnfet$21_15 m1_n1989_16202# m1_n1989_16202# vss vss m1_n2507_16398# vss nfet$21
Xnfet$11_7 m1_32330_25662# m1_32554_23922# m1_32818_24542# vss nfet$11
Xpfet$31_1 vdd m1_n4485_20152# vdd m1_n3206_20274# pfet$31
Xpfet$24_0 vdd vdd m1_n7320_25516# m1_n7186_25858# pfet$24
Xnfet$3_3 m1_9418_21590# m1_9418_21590# m1_9645_21447# m1_9645_21447# m1_9877_21586#
+ vss nfet$3
Xpfet$10_6 vdd vdd m1_32818_24542# m1_33174_24224# pfet$10
Xpfet$5_14 vdd vdd m1_19969_21590# m1_19839_21786# pfet$5
Xnfet$1_0 m1_4509_24346# m1_4509_24346# vss vss m1_3991_24542# vss nfet$1
Xpfet$9_0 vdd vdd m1_n647_25662# m1_n789_25858# pfet$9
Xpfet$2_15 vdd vdd m1_5302_17714# m1_5761_16080# pfet$2
Xpfet$2_26 vdd vdd m1_4832_17714# m1_5302_17714# pfet$2
Xpfet$2_37 vdd m1_7555_16080# m1_7088_18030# m1_6116_17343# pfet$2
Xpfet$2_48 vdd vdd m1_n3064_17714# m1_n2605_16080# pfet$2
Xpfet$2_59 vdd vdd m1_n2605_16080# m1_n7513_20152# pfet$2
Xnfet$29_8 m1_n4623_25487# vss m1_n4464_25980# vss nfet$29
Xpfet$2_7 vdd vdd m1_6275_17836# m1_6116_17343# pfet$2
Xnfet$1_20 m1_21241_24346# m1_21241_24346# m1_20126_25858# m1_20126_25858# m1_22188_25502#
+ vss nfet$1
Xpfet$2_103 vdd m1_14743_16202# m1_14258_17518# m1_14641_17836# pfet$2
Xnfet$21_27 m1_18310_16080# m1_18310_16080# vss vss m1_19873_17358# vss nfet$21
Xnfet$21_16 m1_19747_15778# m1_19747_15778# m1_19637_18030# m1_19637_18030# m1_19873_17358#
+ vss nfet$21
Xnfet$18_1 m1_30256_19792# vss m1_32818_20470# vss nfet$18
Xnfet$5_7 m1_9485_17714# vss m1_10075_17518# vss nfet$5
Xnfet$25_2 m1_n6788_16080# m1_n6788_16080# m1_n7247_17714# m1_n7247_17714# m1_n6690_16398#
+ vss nfet$25
Xpfet$19_3 vdd m1_n5461_18030# vdd m1_n6788_16080# pfet$19
Xpfet$26_4 vdd vdd m1_n4485_21904# m1_n3822_21786# pfet$26
Xpfet$17_0 vdd vdd fout m1_34093_22102# pfet$17
Xpfet$31_2 vdd m1_n5227_20152# vdd m1_n1927_20274# pfet$31
Xnfet$30_0 m1_n9952_24224# m1_n9952_24224# m1_n10308_24542# m1_n10308_24542# m1_n9854_24542#
+ vss nfet$30
Xpfet$24_1 vdd vdd m1_n6111_25858# m1_n6856_24542# pfet$24
Xnfet$3_4 m1_5901_21590# m1_5901_21590# m1_7388_22513# m1_7388_22513# m1_6360_21586#
+ vss nfet$3
Xpfet$10_7 vdd m1_32818_24542# vdd m1_33790_24346# pfet$10
Xpfet$5_15 vdd vdd m1_27003_21590# m1_26873_21786# pfet$5
Xnfet$1_1 m1_3893_24224# m1_3893_24224# m1_3537_24542# m1_3537_24542# m1_3991_24542#
+ vss nfet$1
Xpfet$9_1 vdd vdd m1_n1134_25662# m1_n1271_25858# pfet$9
Xpfet$2_16 vdd vdd m1_3989_15778# m1_1119_17714# pfet$2
Xpfet$2_27 vdd m1_2194_16202# m1_1709_17518# m1_2092_17836# pfet$2
Xpfet$2_38 vdd vdd m1_7088_18030# m1_7198_15778# pfet$2
Xpfet$2_49 vdd m1_n194_15778# m1_n811_16080# m1_n2091_17836# pfet$2
Xpfet$2_8 vdd vdd m1_9331_15478# sd5 pfet$2
Xnfet$29_9 m1_n3184_24224# vss m1_n3541_23922# vss nfet$29
Xnfet$1_21 m1_28991_24224# m1_28991_24224# m1_28635_24542# m1_28635_24542# m1_29089_24542#
+ vss nfet$1
Xnfet$1_10 m1_17546_25658# m1_17546_25658# vss vss m1_18005_25502# vss nfet$1
Xpfet$2_104 vdd vdd m1_14127_16080# m1_n7513_20152# pfet$2
Xnfet$21_17 m1_22493_16080# m1_22493_16080# vss vss m1_24056_17358# vss nfet$21
Xnfet$18_2 m1_31535_19792# m1_32818_20470# vss vss nfet$18
Xpfet$19_4 vdd vdd m1_26217_17714# m1_26676_16080# pfet$19
Xnfet$25_3 m1_n6172_16202# m1_n6172_16202# vss vss m1_n6690_16398# vss nfet$25
Xpfet$26_5 vdd m1_n6839_21786# vdd m1_n5764_21786# pfet$26
Xnfet$5_8 m1_7555_16080# vss m1_7198_15778# vss nfet$5
Xpfet$31_3 vdd m1_n6839_20152# vdd m1_n927_19404# pfet$31
Xnfet$23_0 m1_35837_22102# vss m1_n7513_20152# vss nfet$23
Xnfet$30_1 m1_n9336_24346# m1_n9336_24346# m1_n8625_26174# m1_n8625_26174# m1_n8389_25502#
+ vss nfet$30
Xnfet$3_5 m1_2254_21786# m1_2254_21786# m1_3871_22513# m1_3871_22513# m1_3475_21586#
+ vss nfet$3
Xpfet$5_16 vdd vdd m1_29256_21786# m1_28624_21786# pfet$5
Xnfet$1_2 m1_4997_25658# m1_4997_25658# vss vss m1_5456_25502# vss nfet$1
Xnfet$4_10 m1_9015_17714# m1_9015_17714# vss vss m1_14005_20470# vss nfet$4
Xpfet$9_2 vdd vdd m1_n1271_25858# m1_n10452_25858# pfet$9
Xpfet$2_17 vdd vdd m1_n2091_17836# m1_n2250_17343# pfet$2
Xpfet$2_9 vdd vdd m1_8172_15778# m1_5302_17714# pfet$2
Xpfet$2_28 vdd m1_2905_18030# vdd m1_1578_16080# pfet$2
Xpfet$2_39 vdd m1_7088_18030# vdd m1_5761_16080# pfet$2
Xnfet$1_22 m1_29607_24346# m1_29607_24346# vss vss m1_29089_24542# vss nfet$1
Xnfet$1_11 m1_16442_24224# m1_16442_24224# m1_16086_24542# m1_16086_24542# m1_16540_24542#
+ vss nfet$1
Xpfet$2_105 vdd vdd m1_14258_17518# m1_13668_17714# pfet$2
Xnfet$18_3 m1_30256_22102# vss m1_32818_21586# vss nfet$18
Xnfet$21_18 m1_23930_15778# m1_23930_15778# m1_23820_18030# m1_23820_18030# m1_24056_17358#
+ vss nfet$21
Xnfet$25_4 m1_28113_15778# m1_28113_15778# m1_28003_18030# m1_28003_18030# m1_28239_17358#
+ vss nfet$25
Xpfet$19_5 vdd m1_26217_17714# vdd m1_27292_16202# pfet$19
Xpfet$26_6 vdd vdd m1_n6973_21481# m1_n6839_21786# pfet$26
Xnfet$5_9 sd5 vss m1_9331_15478# vss nfet$5
Xnfet$7_10 m1_26063_15478# vss m1_29239_20152# vss nfet$7
Xnfet$16_0 m1_34843_21786# m1_34843_21786# m1_34093_22102# m1_34093_22102# m1_34329_21430#
+ vss nfet$16
Xpfet$31_4 vdd vdd m1_n6839_20152# m1_n6973_21481# pfet$31
Xnfet$30_2 m1_n8848_25658# m1_n8848_25658# vss vss m1_n8389_25502# vss nfet$30
Xnfet$3_6 m1_2384_21590# m1_2384_21590# m1_3871_22513# m1_3871_22513# m1_2843_21586#
+ vss nfet$3
Xpfet$5_17 vdd vdd m1_25739_21786# m1_25107_21786# pfet$5
Xpfet$22_0 vdd vdd vdd m1_n6624_23622# m1_n7082_23622# m1_n7082_23622# pfet$22
Xnfet$1_3 m1_4509_24346# m1_4509_24346# m1_3394_25858# m1_3394_25858# m1_5456_25502#
+ vss nfet$1
Xnfet$4_11 m1_13198_17714# m1_13198_17714# vss vss m1_17522_20470# vss nfet$4
Xpfet$9_3 vdd vdd m1_1607_24542# m1_n789_25858# pfet$9
Xpfet$2_18 vdd m1_1119_17714# vdd m1_2194_16202# pfet$2
Xpfet$2_29 vdd vdd m1_1578_16080# m1_n7513_20152# pfet$2
Xpfet$7_0 vdd vdd m1_2384_19550# m1_n3534_17714# pfet$7
Xnfet$1_23 m1_25424_24346# m1_25424_24346# m1_24309_25858# m1_24309_25858# m1_26371_25502#
+ vss nfet$1
Xnfet$1_12 m1_17058_24346# m1_17058_24346# m1_15943_25858# m1_15943_25858# m1_18005_25502#
+ vss nfet$1
Xpfet$2_106 vdd vdd m1_14482_17343# m1_17381_17714# pfet$2
Xpfet$19_6 vdd vdd m1_28003_18030# m1_28113_15778# pfet$19
Xnfet$25_5 m1_26676_16080# m1_26676_16080# vss vss m1_28239_17358# vss nfet$25
Xpfet$26_7 vdd vdd m1_n6839_21786# m1_n6380_21786# pfet$26
Xnfet$21_19 m1_23109_16202# m1_23109_16202# vss vss m1_22591_16398# vss nfet$21
Xnfet$16_1 m1_28490_22513# m1_28490_22513# vss vss m1_34329_21430# vss nfet$16
Xnfet$7_11 m1_9331_15478# vss m1_15171_20152# vss nfet$7
Xnfet$30_3 m1_n9336_24346# m1_n9336_24346# vss vss m1_n9854_24542# vss nfet$30
Xnfet$3_7 m1_5771_21786# m1_5771_21786# m1_7388_22513# m1_7388_22513# m1_6992_21586#
+ vss nfet$3
Xpfet$15_0 vdd m1_34093_22102# vdd m1_28490_22513# pfet$15
Xnfet$1_4 m1_12259_24224# m1_12259_24224# m1_11903_24542# m1_11903_24542# m1_12357_24542#
+ vss nfet$1
Xpfet$22_1 vdd m1_n6856_24542# m1_n6856_24542# m1_n6624_23622# m1_n8283_19850# m1_n8283_19850#
+ pfet$22
Xnfet$4_12 m1_16452_19550# m1_16452_19550# vss vss m1_16890_20470# vss nfet$4
Xpfet$9_4 vdd vdd m1_488_21786# m1_n789_25858# pfet$9
Xpfet$2_19 vdd m1_3015_15778# m1_2194_16202# m1_1933_17343# pfet$2
Xpfet$7_1 vdd vdd m1_4620_20152# m1_n3218_15478# pfet$7
Xnfet$1_24 m1_30095_25658# m1_30095_25658# vss vss m1_30554_25502# vss nfet$1
Xnfet$1_13 m1_13363_25658# m1_13363_25658# vss vss m1_13822_25502# vss nfet$1
Xpfet$2_107 vdd m1_15921_16080# m1_15454_18030# m1_14482_17343# pfet$2
Xpfet$19_7 vdd m1_28003_18030# vdd m1_26676_16080# pfet$19
Xnfet$25_6 m1_27292_16202# m1_27292_16202# vss vss m1_26774_16398# vss nfet$25
Xnfet$16_2 m1_9645_21447# m1_9645_21447# vss vss m1_30492_21430# vss nfet$16
Xnfet$7_12 m1_13514_15478# vss m1_18688_20152# vss nfet$7
Xnfet$30_4 m1_n4978_24224# m1_n4978_24224# m1_n10452_25858# m1_n10452_25858# m1_n4880_24542#
+ vss nfet$30
Xnfet$3_8 m1_23486_21590# m1_23486_21590# m1_24973_22513# m1_24973_22513# m1_23945_21586#
+ vss nfet$3
Xpfet$15_1 vdd vdd m1_34093_22102# m1_34843_21786# pfet$15
Xnfet$1_5 m1_8692_24346# m1_8692_24346# vss vss m1_8174_24542# vss nfet$1
Xnfet$21_0 m1_7198_15778# m1_7198_15778# m1_7088_18030# m1_7088_18030# m1_7324_17358#
+ vss nfet$21
Xnfet$4_13 m1_19969_19550# m1_19969_19550# vss vss m1_20407_20470# vss nfet$4
Xpfet$9_5 vdd vdd m1_326_24346# m1_n7513_20152# pfet$9
Xpfet$7_2 vdd vdd m1_1103_20152# m1_n7401_15478# pfet$7
Xnfet$1_25 m1_29607_24346# m1_29607_24346# m1_28492_25858# m1_28492_25858# m1_30554_25502#
+ vss nfet$1
Xnfet$1_14 m1_12875_24346# m1_12875_24346# m1_11760_25858# m1_11760_25858# m1_13822_25502#
+ vss nfet$1
Xpfet$3_30 vdd vdd vdd m1_17539_22402# m1_16322_21786# m1_16322_21786# pfet$3
Xpfet$2_108 vdd vdd m1_15454_18030# m1_15564_15778# pfet$2
Xnfet$25_7 m1_26676_16080# m1_26676_16080# m1_26217_17714# m1_26217_17714# m1_26774_16398#
+ vss nfet$25
Xnfet$7_13 m1_13198_17714# vss m1_16452_19550# vss nfet$7
Xnfet$30_5 m1_n4362_24346# m1_n4362_24346# vss vss m1_n4880_24542# vss nfet$30
Xnfet$16_3 m1_7388_22513# m1_7388_22513# m1_30256_22102# m1_30256_22102# m1_30492_21430#
+ vss nfet$16
Xnfet$3_9 m1_23356_21786# m1_23356_21786# m1_24973_22513# m1_24973_22513# m1_24577_21586#
+ vss nfet$3
Xpfet$15_2 vdd vdd m1_30256_22102# m1_7388_22513# pfet$15
Xnfet$21_1 m1_5761_16080# m1_5761_16080# vss vss m1_7324_17358# vss nfet$21
Xnfet$14_0 m1_11039_21786# m1_11039_21786# vss vss m1_9877_21586# vss nfet$14
Xnfet$1_6 m1_8076_24224# m1_8076_24224# m1_7720_24542# m1_7720_24542# m1_8174_24542#
+ vss nfet$1
Xnfet$4_14 m1_17381_17714# m1_17381_17714# vss vss m1_21039_20470# vss nfet$4
Xpfet$9_6 vdd vdd m1_n290_24224# m1_n910_23922# pfet$9
Xpfet$20_0 vdd m1_n4377_15778# m1_n4994_16080# m1_n6274_17836# pfet$20
Xnfet$14_10 m1_21590_21786# m1_21590_21786# vss vss m1_20428_21586# vss nfet$14
Xpfet$7_3 vdd vdd m1_5901_19550# m1_649_17714# pfet$7
Xnfet$1_26 m1_25912_25658# m1_25912_25658# vss vss m1_26371_25502# vss nfet$1
Xnfet$1_15 m1_25424_24346# m1_25424_24346# vss vss m1_24906_24542# vss nfet$1
Xpfet$3_31 vdd vdd vdd m1_27462_22102# m1_27003_21590# m1_27003_21590# pfet$3
Xpfet$3_20 vdd vdd vdd m1_20428_22102# m1_19969_21590# m1_19969_21590# pfet$3
Xpfet$2_109 vdd vdd m1_10299_17343# m1_13198_17714# pfet$2
Xpfet$5_0 vdd vdd m1_n1133_21590# m1_n1263_21786# pfet$5
Xnfet$2_80 m1_28147_25662# m1_28991_24224# m1_30095_25658# vss nfet$2
Xnfet$7_14 m1_21564_17714# vss m1_23486_19550# vss nfet$7
Xnfet$30_6 m1_n4978_24224# m1_n4978_24224# vss vss m1_n3415_25502# vss nfet$30
Xnfet$22_10 m1_9331_15478# m1_9331_15478# m1_n3822_21786# m1_n3822_21786# m1_13373_20470#
+ vss nfet$22
Xnfet$8_0 sd9 vss m1_n7401_15478# vss nfet$8
Xpfet$15_3 vdd m1_31535_22102# vdd m1_3871_22513# pfet$15
Xnfet$21_2 m1_9944_16080# m1_9944_16080# vss vss m1_11507_17358# vss nfet$21
Xnfet$14_1 m1_11671_21786# m1_11671_21786# vss vss m1_10509_21586# vss nfet$14
Xnfet$1_7 m1_9180_25658# m1_9180_25658# vss vss m1_9639_25502# vss nfet$1
Xnfet$4_15 m1_21564_17714# m1_21564_17714# vss vss m1_24556_20470# vss nfet$4
Xpfet$9_7 vdd vdd m1_32330_25662# m1_32193_25858# pfet$9
Xpfet$20_1 vdd m1_n5351_15778# m1_n6172_16202# m1_n6433_17343# pfet$20
Xpfet$13_0 vdd m1_n647_25662# m1_n910_23922# m1_n1134_25662# pfet$13
Xpfet$7_4 vdd vdd m1_12935_19550# m1_9015_17714# pfet$7
Xnfet$14_11 m1_22222_21786# m1_22222_21786# vss vss m1_21060_21586# vss nfet$14
Xnfet$5_80 m1_18824_17836# m1_19747_15778# m1_18926_16202# vss nfet$5
Xnfet$1_27 m1_12875_24346# m1_12875_24346# vss vss m1_12357_24542# vss nfet$1
Xpfet$3_32 vdd m1_28490_22513# m1_28490_22513# m1_28090_22402# m1_28624_21786# m1_28624_21786#
+ pfet$3
Xnfet$1_16 m1_24808_24224# m1_24808_24224# m1_24452_24542# m1_24452_24542# m1_24906_24542#
+ vss nfet$1
Xpfet$3_21 vdd vdd vdd m1_21056_22402# m1_19839_21786# m1_19839_21786# pfet$3
Xpfet$3_10 vdd m1_3871_22513# m1_3871_22513# m1_2843_22102# m1_4637_21786# m1_4637_21786#
+ pfet$3
Xpfet$5_1 vdd vdd m1_11671_21786# m1_11039_21786# pfet$5
Xpfet$1_110 vdd m1_11903_24542# vdd m1_12875_24346# pfet$1
Xnfet$2_81 m1_n7513_20152# vss m1_25424_24346# vss nfet$2
Xnfet$2_70 m1_21590_21786# vss m1_28010_25858# vss nfet$2
Xnfet$37_0 m1_n6839_20152# vss m1_n8145_21908# vss nfet$37
Xnfet$7_15 m1_17697_15478# vss m1_22205_20152# vss nfet$7
Xnfet$30_7 m1_n3541_23922# m1_n3541_23922# m1_n3651_26174# m1_n3651_26174# m1_n3415_25502#
+ vss nfet$30
Xnfet$22_11 m1_15171_20152# m1_15171_20152# m1_n3822_21786# m1_n3822_21786# m1_14005_20470#
+ vss nfet$22
Xnfet$8_1 sd2 vss m1_21880_15478# vss nfet$8
Xpfet$15_4 vdd m1_30256_22102# vdd m1_9645_21447# pfet$15
Xnfet$1_8 m1_8692_24346# m1_8692_24346# m1_7577_25858# m1_7577_25858# m1_9639_25502#
+ vss nfet$1
Xnfet$21_3 m1_11381_15778# m1_11381_15778# m1_11271_18030# m1_11271_18030# m1_11507_17358#
+ vss nfet$21
Xnfet$14_2 m1_8154_21786# m1_8154_21786# vss vss m1_6992_21586# vss nfet$14
Xnfet$4_16 m1_23486_19550# m1_23486_19550# vss vss m1_23924_20470# vss nfet$4
Xpfet$9_8 vdd vdd m1_33174_24224# m1_32554_23922# pfet$9
Xpfet$6_10 vdd vdd m1_27031_17343# m1_n10452_25858# pfet$6
Xpfet$20_2 vdd m1_n4994_16080# m1_n5461_18030# m1_n6433_17343# pfet$20
Xpfet$13_1 vdd m1_n910_23922# m1_n646_24542# m1_n1271_25858# pfet$13
Xpfet$7_5 vdd vdd m1_8137_20152# m1_965_15478# pfet$7
Xnfet$5_81 m1_13198_17714# vss m1_10299_17343# vss nfet$5
Xnfet$14_12 m1_18073_21786# m1_18073_21786# vss vss m1_16911_21586# vss nfet$14
Xnfet$5_70 m1_n7513_20152# vss m1_18310_16080# vss nfet$5
Xpfet$3_33 vdd m1_28490_22513# m1_28490_22513# m1_27462_22102# m1_29256_21786# m1_29256_21786#
+ pfet$3
Xnfet$1_17 m1_20625_24224# m1_20625_24224# m1_20269_24542# m1_20269_24542# m1_20723_24542#
+ vss nfet$1
Xpfet$3_22 vdd m1_21456_22513# m1_21456_22513# m1_20428_22102# m1_22222_21786# m1_22222_21786#
+ pfet$3
Xpfet$3_11 vdd vdd vdd m1_2843_22102# m1_2384_21590# m1_2384_21590# pfet$3
Xpfet$5_2 vdd vdd m1_12935_21590# m1_12805_21786# pfet$5
Xpfet$1_100 vdd vdd m1_29607_24346# m1_n7513_20152# pfet$1
Xnfet$2_82 m1_11415_25662# m1_12259_24224# m1_13363_25658# vss nfet$2
Xnfet$2_71 m1_28147_25662# m1_28371_23922# m1_28635_24542# vss nfet$2
Xnfet$2_60 pd6 vss m1_16322_21786# vss nfet$2
Xpfet$9_10 vdd vdd m1_35071_24542# m1_32675_25947# pfet$9
Xnfet$7_16 m1_17381_17714# vss m1_19969_19550# vss nfet$7
Xnfet$8_2 sd1 vss m1_26063_15478# vss nfet$8
Xnfet$22_12 m1_18688_20152# m1_18688_20152# m1_n1927_20274# m1_n1927_20274# m1_17522_20470#
+ vss nfet$22
Xnfet$1_9 m1_17058_24346# m1_17058_24346# vss vss m1_16540_24542# vss nfet$1
Xnfet$21_4 m1_10560_16202# m1_10560_16202# vss vss m1_10042_16398# vss nfet$21
Xnfet$14_3 m1_7522_21786# m1_7522_21786# vss vss m1_6360_21586# vss nfet$14
Xnfet$4_17 m1_12935_19550# m1_12935_19550# vss vss m1_13373_20470# vss nfet$4
Xpfet$9_9 vdd vdd m1_28624_21786# m1_32675_25947# pfet$9
Xpfet$6_11 vdd vdd m1_26807_17518# m1_26217_17714# pfet$6
Xnfet$12_0 pd1 vss m1_n1263_21786# vss nfet$12
Xpfet$20_3 vdd m1_n6172_16202# m1_n6657_17518# m1_n6274_17836# pfet$20
Xpfet$13_2 vdd m1_n290_24224# m1_814_25658# m1_n1271_25858# pfet$13
Xnfet$5_82 m1_10299_17343# vss m1_10458_17836# vss nfet$5
Xnfet$14_13 m1_18705_21786# m1_18705_21786# vss vss m1_17543_21586# vss nfet$14
Xnfet$5_71 m1_14641_17836# m1_15921_16080# m1_15454_18030# vss nfet$5
Xnfet$5_60 m1_18665_17343# vss m1_18824_17836# vss nfet$5
Xpfet$7_6 vdd vdd m1_9418_19550# m1_4832_17714# pfet$7
Xnfet$1_18 m1_21241_24346# m1_21241_24346# vss vss m1_20723_24542# vss nfet$1
Xpfet$3_12 vdd vdd vdd m1_3471_22402# m1_2254_21786# m1_2254_21786# pfet$3
Xpfet$3_34 vdd vdd vdd m1_28090_22402# m1_26873_21786# m1_26873_21786# pfet$3
Xpfet$3_23 vdd vdd vdd m1_23945_22102# m1_23486_21590# m1_23486_21590# pfet$3
Xpfet$5_3 vdd vdd m1_9418_21590# m1_9288_21786# pfet$5
Xpfet$1_101 vdd vdd m1_28010_25858# m1_21590_21786# pfet$1
Xnfet$2_72 m1_23827_25858# m1_25912_25658# m1_26705_24542# vss nfet$2
Xnfet$2_61 m1_23964_25662# m1_24808_24224# m1_25912_25658# vss nfet$2
Xnfet$2_50 m1_n7513_20152# vss m1_21241_24346# vss nfet$2
Xpfet$3_0 vdd vdd vdd m1_n674_22102# m1_n1133_21590# m1_n1133_21590# pfet$3
Xnfet$7_17 m1_21880_15478# vss m1_25722_20152# vss nfet$7
Xpfet$9_11 vdd vdd m1_32817_25662# m1_32675_25947# pfet$9
Xnfet$22_13 m1_13514_15478# m1_13514_15478# m1_n1927_20274# m1_n1927_20274# m1_16890_20470#
+ vss nfet$22
Xpfet$29_0 vdd vdd vdd m1_n8047_19550# m1_n7513_20152# m1_n7513_20152# pfet$29
Xnfet$21_5 m1_9944_16080# m1_9944_16080# m1_9485_17714# m1_9485_17714# m1_10042_16398#
+ vss nfet$21
Xnfet$14_4 m1_1120_21786# m1_1120_21786# vss vss m1_n42_21586# vss nfet$14
Xnfet$6_0 m1_n1263_21786# vss m1_n1133_21590# vss nfet$6
Xpfet$6_12 vdd vdd m1_26676_16080# m1_n7513_20152# pfet$6
Xpfet$20_4 vdd m1_28113_15778# m1_27292_16202# m1_27031_17343# pfet$20
Xpfet$13_3 vdd m1_814_25658# m1_1607_24542# m1_n1134_25662# pfet$13
Xnfet$12_1 pd2 vss m1_2254_21786# vss nfet$12
Xpfet$11_0 vdd vdd vdd m1_33050_22344# m1_31535_22102# m1_31535_22102# pfet$11
Xnfet$14_14 m1_15188_21786# m1_15188_21786# vss vss m1_14026_21586# vss nfet$14
Xnfet$5_72 m1_17851_17714# vss m1_18441_17518# vss nfet$5
Xnfet$5_61 m1_20104_16080# vss m1_19747_15778# vss nfet$5
Xnfet$5_50 m1_25747_17714# vss m1_22848_17343# vss nfet$5
Xpfet$7_7 vdd vdd m1_11654_20152# m1_5148_15478# pfet$7
Xnfet$1_19 m1_21729_25658# m1_21729_25658# vss vss m1_22188_25502# vss nfet$1
Xpfet$27_10 vdd vdd m1_n10933_25858# fin pfet$27
Xpfet$3_35 vdd vdd vdd m1_13394_22102# m1_12935_21590# m1_12935_21590# pfet$3
Xpfet$3_24 vdd m1_17939_22513# m1_17939_22513# m1_16911_22102# m1_18705_21786# m1_18705_21786#
+ pfet$3
Xpfet$3_13 vdd vdd vdd m1_6988_22402# m1_5771_21786# m1_5771_21786# pfet$3
Xpfet$5_4 vdd vdd m1_8154_21786# m1_7522_21786# pfet$5
Xpfet$1_102 vdd m1_28371_23922# m1_28635_24542# m1_28010_25858# pfet$1
Xnfet$2_73 m1_24309_25858# vss m1_21590_21786# vss nfet$2
Xnfet$2_62 m1_24188_23922# vss m1_24808_24224# vss nfet$2
Xnfet$2_51 m1_19644_25858# m1_21729_25658# m1_22522_24542# vss nfet$2
Xnfet$2_40 m1_15598_25662# m1_16442_24224# m1_17546_25658# vss nfet$2
Xpfet$3_1 vdd m1_7388_22513# m1_7388_22513# m1_6988_22402# m1_7522_21786# m1_7522_21786#
+ pfet$3
Xpfet$9_12 vdd vdd m1_32193_25858# m1_25107_21786# pfet$9
Xnfet$22_14 m1_22205_20152# m1_22205_20152# m1_n2543_20130# m1_n2543_20130# m1_21039_20470#
+ vss nfet$22
Xpfet$29_1 vdd m1_n8283_19850# m1_n8283_19850# m1_n8047_19550# m1_n8283_20611# m1_n8283_20611#
+ pfet$29
Xnfet$35_0 m1_n927_19404# m1_n927_19404# vss vss m1_n6282_20470# vss nfet$35
Xnfet$21_6 m1_1578_16080# m1_1578_16080# vss vss m1_3141_17358# vss nfet$21
Xnfet$14_5 m1_4005_21786# m1_4005_21786# vss vss m1_2843_21586# vss nfet$14
Xpfet$1_90 vdd vdd m1_24309_25858# m1_25424_24346# pfet$1
Xpfet$6_13 vdd vdd m1_25747_17714# m1_26217_17714# pfet$6
Xnfet$6_1 m1_11039_21786# vss m1_11671_21786# vss nfet$6
Xnfet$12_2 pd9 vss m1_26873_21786# vss nfet$12
Xpfet$13_4 vdd m1_33174_24224# m1_34278_25658# m1_32193_25858# pfet$13
Xpfet$20_5 vdd m1_29087_15778# m1_28470_16080# m1_27190_17836# pfet$20
Xnfet$14_15 m1_14556_21786# m1_14556_21786# vss vss m1_13394_21586# vss nfet$14
Xnfet$5_73 m1_13668_17714# vss m1_16538_15778# vss nfet$5
Xnfet$5_62 m1_18665_17343# m1_20721_15778# m1_20104_16080# vss nfet$5
Xnfet$5_51 m1_n7513_20152# vss m1_22493_16080# vss nfet$5
Xnfet$5_40 m1_n2250_17343# m1_n194_15778# m1_n811_16080# vss nfet$5
Xpfet$7_8 vdd vdd m1_n1133_19550# m1_n7383_17599# pfet$7
Xpfet$3_25 vdd m1_17939_22513# m1_17939_22513# m1_17539_22402# m1_18073_21786# m1_18073_21786#
+ pfet$3
Xpfet$3_14 vdd vdd vdd m1_n46_22402# m1_n1263_21786# m1_n1263_21786# pfet$3
Xpfet$27_11 vdd vdd m1_n9336_24346# vss pfet$27
Xpfet$5_5 vdd vdd m1_1120_21786# m1_488_21786# pfet$5
Xpfet$1_103 vdd vdd m1_28635_24542# m1_28991_24224# pfet$1
Xnfet$2_74 pd8 vss m1_23356_21786# vss nfet$2
Xnfet$2_63 m1_14556_21786# vss m1_19644_25858# vss nfet$2
Xnfet$2_52 m1_20126_25858# vss m1_22522_24542# vss nfet$2
Xnfet$2_41 pd5 vss m1_12805_21786# vss nfet$2
Xnfet$2_30 m1_n7513_20152# vss m1_17058_24346# vss nfet$2
Xpfet$3_2 vdd m1_7388_22513# m1_7388_22513# m1_6360_22102# m1_8154_21786# m1_8154_21786#
+ pfet$3
Xpfet$9_13 vdd vdd m1_33790_24346# m1_n7513_20152# pfet$9
Xnfet$35_1 m1_n2543_20130# m1_n2543_20130# m1_n5227_20152# m1_n5227_20152# m1_n2445_20470#
+ vss nfet$35
Xpfet$29_2 vdd m1_n8283_20611# m1_n8283_20611# m1_n8047_22344# m1_n8145_21908# m1_n8145_21908#
+ pfet$29
Xnfet$22_15 m1_17697_15478# m1_17697_15478# m1_n2543_20130# m1_n2543_20130# m1_20407_20470#
+ vss nfet$22
Xnfet$28_0 m1_n3822_20130# m1_n3822_20130# m1_n4485_20152# m1_n4485_20152# m1_n3724_20470#
+ vss nfet$28
Xnfet$21_7 m1_5761_16080# m1_5761_16080# m1_5302_17714# m1_5302_17714# m1_5859_16398#
+ vss nfet$21
Xnfet$14_6 m1_4637_21786# m1_4637_21786# vss vss m1_3475_21586# vss nfet$14
Xpfet$1_91 vdd vdd m1_23356_21786# pd8 pfet$1
Xpfet$1_80 vdd vdd m1_17058_24346# m1_n7513_20152# pfet$1
Xnfet$6_2 m1_12805_21786# vss m1_12935_21590# vss nfet$6
Xpfet$13_5 vdd m1_32817_25662# m1_32554_23922# m1_32330_25662# pfet$13
Xpfet$20_6 vdd m1_28470_16080# m1_28003_18030# m1_27031_17343# pfet$20
Xnfet$5_74 m1_14482_17343# vss m1_14641_17836# vss nfet$5
Xnfet$5_63 m1_13668_17714# vss m1_14258_17518# vss nfet$5
Xnfet$5_52 m1_23007_17836# m1_24287_16080# m1_23820_18030# vss nfet$5
Xpfet$7_9 vdd vdd m1_27003_19550# m1_25747_17714# pfet$7
Xnfet$5_30 sd6 vss m1_5148_15478# vss nfet$5
Xnfet$5_41 m1_n2091_17836# m1_n1168_15778# m1_n1989_16202# vss nfet$5
Xnfet$14_16 m1_28624_21786# m1_28624_21786# vss vss m1_27462_21586# vss nfet$14
Xnfet$10_0 m1_n10452_25858# vss m1_n1271_25858# vss nfet$10
Xpfet$3_26 vdd vdd vdd m1_16911_22102# m1_16452_21590# m1_16452_21590# pfet$3
Xpfet$3_15 vdd m1_354_22513# m1_354_22513# m1_n46_22402# m1_488_21786# m1_488_21786#
+ pfet$3
Xpfet$27_12 vdd vdd m1_n7082_23622# m1_n8625_26174# pfet$27
Xpfet$5_6 vdd vdd m1_5901_21590# m1_5771_21786# pfet$5
Xpfet$1_104 vdd m1_25912_25658# m1_26705_24542# m1_23964_25662# pfet$1
Xnfet$2_75 m1_28371_23922# vss m1_28991_24224# vss nfet$2
Xnfet$2_64 m1_19644_25858# vss m1_19781_25662# vss nfet$2
Xnfet$2_53 m1_23827_25858# m1_24451_25662# m1_24188_23922# vss nfet$2
Xnfet$2_42 m1_15943_25858# vss m1_16085_25662# vss nfet$2
Xnfet$2_31 m1_15943_25858# vss m1_18339_24542# vss nfet$2
Xnfet$2_20 pd3 vss m1_5771_21786# vss nfet$2
Xpfet$3_3 vdd m1_9645_21447# m1_9645_21447# m1_10505_22402# m1_11039_21786# m1_11039_21786#
+ pfet$3
Xnfet$22_16 m1_25722_20152# m1_25722_20152# m1_n3206_20274# m1_n3206_20274# m1_24556_20470#
+ vss nfet$22
Xnfet$28_1 m1_n1927_20274# m1_n1927_20274# vss vss m1_n2445_20470# vss nfet$28
Xpfet$29_3 vdd vdd vdd m1_n8047_22344# m1_n8283_19850# m1_n8283_19850# pfet$29
Xpfet$1_0 vdd vdd m1_3049_25662# m1_2912_25858# pfet$1
Xpfet$1_92 vdd vdd m1_28492_25858# m1_29607_24346# pfet$1
Xpfet$1_81 vdd vdd m1_18339_24542# m1_15943_25858# pfet$1
Xpfet$1_70 vdd vdd m1_14156_24542# m1_11760_25858# pfet$1
Xnfet$14_7 m1_488_21786# m1_488_21786# vss vss m1_n674_21586# vss nfet$14
Xnfet$21_8 m1_3015_15778# m1_3015_15778# m1_2905_18030# m1_2905_18030# m1_3141_17358#
+ vss nfet$21
Xpfet$27_0 vdd vdd m1_n10796_25662# m1_n10933_25858# pfet$27
Xnfet$6_3 m1_9288_21786# vss m1_9418_21590# vss nfet$6
Xpfet$13_6 vdd m1_34278_25658# m1_35071_24542# m1_32330_25662# pfet$13
Xpfet$20_7 vdd m1_27292_16202# m1_26807_17518# m1_27190_17836# pfet$20
Xnfet$4_0 m1_n3534_17714# m1_n3534_17714# vss vss m1_3454_20470# vss nfet$4
Xnfet$14_17 m1_29256_21786# m1_29256_21786# vss vss m1_28094_21586# vss nfet$14
Xnfet$5_75 sd3 vss m1_17697_15478# vss nfet$5
Xnfet$5_64 m1_13668_17714# vss m1_13198_17714# vss nfet$5
Xnfet$5_53 m1_22848_17343# vss m1_23007_17836# vss nfet$5
Xnfet$5_31 m1_1933_17343# m1_3989_15778# m1_3372_16080# vss nfet$5
Xnfet$5_20 m1_1119_17714# vss m1_1709_17518# vss nfet$5
Xnfet$5_42 m1_n811_16080# vss m1_n1168_15778# vss nfet$5
Xnfet$10_1 m1_n789_25858# vss m1_n647_25662# vss nfet$10
Xpfet$3_27 vdd m1_14422_22513# m1_14422_22513# m1_14022_22402# m1_14556_21786# m1_14556_21786#
+ pfet$3
Xpfet$3_16 vdd m1_24973_22513# m1_24973_22513# m1_23945_22102# m1_25739_21786# m1_25739_21786#
+ pfet$3
Xpfet$27_13 vdd vdd m1_n8055_24542# m1_n8625_26174# pfet$27
Xpfet$5_7 vdd vdd m1_4637_21786# m1_4005_21786# pfet$5
Xpfet$1_105 vdd vdd m1_30888_24542# m1_28492_25858# pfet$1
Xnfet$2_76 m1_28492_25858# vss m1_28634_25662# vss nfet$2
Xnfet$2_65 m1_28492_25858# vss m1_25107_21786# vss nfet$2
Xnfet$2_54 m1_24309_25858# vss m1_24451_25662# vss nfet$2
Xnfet$2_43 m1_15461_25858# vss m1_15598_25662# vss nfet$2
Xnfet$2_32 m1_15461_25858# m1_17546_25658# m1_18339_24542# vss nfet$2
Xnfet$2_21 m1_11278_25858# m1_11902_25662# m1_11639_23922# vss nfet$2
Xnfet$2_10 m1_7577_25858# vss m1_9973_24542# vss nfet$2
Xpfet$3_4 vdd vdd vdd m1_9877_22102# m1_9418_21590# m1_9418_21590# pfet$3
Xnfet$22_17 m1_21880_15478# m1_21880_15478# m1_n3206_20274# m1_n3206_20274# m1_23924_20470#
+ vss nfet$22
Xpfet$1_1 vdd m1_3536_25662# m1_3273_23922# m1_3049_25662# pfet$1
Xnfet$28_2 m1_n3206_20274# m1_n3206_20274# vss vss m1_n3724_20470# vss nfet$28
Xnfet$14_8 m1_25739_21786# m1_25739_21786# vss vss m1_24577_21586# vss nfet$14
Xnfet$21_9 m1_2194_16202# m1_2194_16202# vss vss m1_1676_16398# vss nfet$21
Xpfet$27_1 vdd vdd m1_n10309_25662# m1_n10452_25858# pfet$27
Xpfet$1_93 vdd m1_28991_24224# m1_30095_25658# m1_28010_25858# pfet$1
Xpfet$1_82 vdd vdd m1_21241_24346# m1_n7513_20152# pfet$1
Xpfet$1_71 vdd vdd m1_11039_21786# m1_11760_25858# pfet$1
Xpfet$1_60 vdd vdd m1_20126_25858# m1_21241_24346# pfet$1
Xnfet$33_0 m1_n8283_20611# vss m1_n8283_19850# vss nfet$33
Xnfet$6_4 m1_7522_21786# vss m1_8154_21786# vss nfet$6
Xpfet$13_7 vdd m1_32554_23922# m1_32818_24542# m1_32193_25858# pfet$13
Xnfet$4_1 m1_2384_19550# m1_2384_19550# vss vss m1_2822_20470# vss nfet$4
Xnfet$5_76 m1_14482_17343# m1_16538_15778# m1_15921_16080# vss nfet$5
Xnfet$5_65 m1_14482_17343# m1_14743_16202# m1_14258_17518# vss nfet$5
Xnfet$5_54 m1_22848_17343# m1_23109_16202# m1_22624_17518# vss nfet$5
Xnfet$5_32 m1_2092_17836# m1_3015_15778# m1_2194_16202# vss nfet$5
Xnfet$5_21 m1_1933_17343# m1_2194_16202# m1_1709_17518# vss nfet$5
Xnfet$5_10 m1_11738_16080# vss m1_11381_15778# vss nfet$5
Xnfet$5_43 sd8 vss m1_n3218_15478# vss nfet$5
Xnfet$10_2 m1_n1271_25858# vss m1_n1134_25662# vss nfet$10
Xpfet$3_28 vdd m1_14422_22513# m1_14422_22513# m1_13394_22102# m1_15188_21786# m1_15188_21786#
+ pfet$3
Xpfet$3_17 vdd m1_21456_22513# m1_21456_22513# m1_21056_22402# m1_21590_21786# m1_21590_21786#
+ pfet$3
Xpfet$5_8 vdd vdd m1_2384_21590# m1_2254_21786# pfet$5
Xpfet$1_106 vdd vdd m1_25107_21786# m1_28492_25858# pfet$1
Xnfet$2_44 m1_15822_23922# vss m1_16442_24224# vss nfet$2
Xnfet$2_33 m1_11760_25858# vss m1_14156_24542# vss nfet$2
Xnfet$2_22 m1_11760_25858# vss m1_11902_25662# vss nfet$2
Xnfet$2_11 m1_7522_21786# vss m1_11278_25858# vss nfet$2
Xnfet$2_77 m1_28010_25858# vss m1_28147_25662# vss nfet$2
Xnfet$2_66 m1_28010_25858# m1_30095_25658# m1_30888_24542# vss nfet$2
Xnfet$2_55 m1_23827_25858# vss m1_23964_25662# vss nfet$2
Xpfet$3_5 vdd m1_9645_21447# m1_9645_21447# m1_9877_22102# m1_11671_21786# m1_11671_21786#
+ pfet$3
Xnfet$28_3 m1_n6973_21481# m1_n6973_21481# m1_n6839_20152# m1_n6839_20152# m1_n6282_20470#
+ vss nfet$28
Xpfet$1_2 vdd vdd m1_3394_25858# m1_4509_24346# pfet$1
Xnfet$14_9 m1_25107_21786# m1_25107_21786# vss vss m1_23945_21586# vss nfet$14
Xpfet$1_94 vdd m1_28492_25858# vdd m1_30095_25658# pfet$1
Xpfet$1_83 vdd m1_21729_25658# m1_22522_24542# m1_19781_25662# pfet$1
Xpfet$1_72 vdd m1_13363_25658# m1_14156_24542# m1_11415_25662# pfet$1
Xpfet$1_61 vdd m1_24452_24542# vdd m1_25424_24346# pfet$1
Xpfet$1_50 vdd vdd m1_20268_25662# m1_20126_25858# pfet$1
Xnfet$33_1 m1_n7513_20152# m1_n8283_19850# vss vss nfet$33
Xnfet$26_0 m1_n10452_25858# m1_n10452_25858# m1_n7186_25858# m1_n7186_25858# m1_n6629_25502#
+ vss nfet$26
Xpfet$27_2 vdd vdd m1_n9952_24224# m1_n10572_23922# pfet$27
Xnfet$6_5 m1_488_21786# vss m1_1120_21786# vss nfet$6
Xpfet$32_0 vdd vdd vdd m1_n5019_19550# m1_n4485_20152# m1_n4485_20152# pfet$32
Xnfet$4_2 m1_5901_19550# m1_5901_19550# vss vss m1_6339_20470# vss nfet$4
Xnfet$5_77 sd4 vss m1_13514_15478# vss nfet$5
Xnfet$5_66 m1_n7513_20152# vss m1_14127_16080# vss nfet$5
Xnfet$5_55 m1_22034_17714# vss m1_24904_15778# vss nfet$5
Xnfet$5_44 m1_n2091_17836# m1_n811_16080# m1_n1278_18030# vss nfet$5
Xnfet$5_33 sd7 vss m1_965_15478# vss nfet$5
Xnfet$5_22 m1_6116_17343# m1_6377_16202# m1_5892_17518# vss nfet$5
Xnfet$5_11 m1_10299_17343# m1_12355_15778# m1_11738_16080# vss nfet$5
Xnfet$10_3 m1_n7513_20152# vss m1_326_24346# vss nfet$10
Xpfet$3_29 vdd vdd vdd m1_14022_22402# m1_12805_21786# m1_12805_21786# pfet$3
Xpfet$5_9 vdd vdd m1_22222_21786# m1_21590_21786# pfet$5
Xpfet$3_18 vdd vdd vdd m1_24573_22402# m1_23356_21786# m1_23356_21786# pfet$3
Xpfet$1_107 vdd m1_24309_25858# vdd m1_25912_25658# pfet$1
Xnfet$2_78 m1_28010_25858# m1_28634_25662# m1_28371_23922# vss nfet$2
Xnfet$2_67 m1_28492_25858# vss m1_30888_24542# vss nfet$2
Xnfet$2_56 m1_19781_25662# m1_20625_24224# m1_21729_25658# vss nfet$2
Xnfet$2_45 m1_15461_25858# m1_16085_25662# m1_15822_23922# vss nfet$2
Xnfet$2_34 m1_11278_25858# m1_13363_25658# m1_14156_24542# vss nfet$2
Xnfet$2_23 m1_11278_25858# vss m1_11415_25662# vss nfet$2
Xnfet$2_12 m1_7577_25858# vss m1_7522_21786# vss nfet$2
Xpfet$3_6 vdd vdd vdd m1_10505_22402# m1_9288_21786# m1_9288_21786# pfet$3
Xnfet$28_4 m1_2590_19404# m1_2590_19404# vss vss m1_n2445_21430# vss nfet$28
Xpfet$1_3 vdd m1_3394_25858# vdd m1_4997_25658# pfet$1
Xpfet$1_95 vdd vdd m1_28991_24224# m1_28371_23922# pfet$1
Xnfet$19_0 m1_34093_22102# vss fout vss nfet$19
Xpfet$1_84 vdd vdd m1_23827_25858# m1_18073_21786# pfet$1
Xpfet$1_73 vdd m1_16086_24542# vdd m1_17058_24346# pfet$1
Xpfet$1_62 vdd vdd m1_24452_24542# m1_24808_24224# pfet$1
Xpfet$1_51 vdd vdd m1_20625_24224# m1_20005_23922# pfet$1
Xpfet$1_40 vdd vdd m1_11760_25858# m1_12875_24346# pfet$1
Xnfet$33_2 m1_n8145_21908# vss m1_n8283_20611# vss nfet$33
Xpfet$27_3 vdd vdd m1_n4978_24224# vss pfet$27
Xnfet$26_1 m1_n6111_25858# m1_n6111_25858# vss vss m1_n6629_25502# vss nfet$26
Xnfet$6_6 m1_5771_21786# vss m1_5901_21590# vss nfet$6
Xpfet$25_0 vdd vdd m1_n8625_26174# m1_n9336_24346# pfet$25
Xnfet$4_3 m1_4832_17714# m1_4832_17714# vss vss m1_10488_20470# vss nfet$4
Xnfet$5_78 m1_14641_17836# m1_15564_15778# m1_14743_16202# vss nfet$5
Xnfet$5_67 m1_17381_17714# vss m1_14482_17343# vss nfet$5
Xnfet$5_56 m1_24287_16080# vss m1_23930_15778# vss nfet$5
Xnfet$5_45 m1_n3064_17714# vss m1_n194_15778# vss nfet$5
Xnfet$5_34 m1_n2250_17343# vss m1_n2091_17836# vss nfet$5
Xnfet$5_23 m1_5302_17714# vss m1_4832_17714# vss nfet$5
Xnfet$5_12 m1_9485_17714# vss m1_12355_15778# vss nfet$5
Xnfet$10_4 m1_n789_25858# vss m1_1607_24542# vss nfet$10
Xpfet$3_19 vdd m1_24973_22513# m1_24973_22513# m1_24573_22402# m1_25107_21786# m1_25107_21786#
+ pfet$3
Xnfet$2_0 m1_3394_25858# vss m1_5790_24542# vss nfet$2
Xpfet$1_108 vdd vdd m1_25424_24346# m1_n7513_20152# pfet$1
Xnfet$2_79 pd7 vss m1_19839_21786# vss nfet$2
Xnfet$2_68 m1_n7513_20152# vss m1_29607_24346# vss nfet$2
Xnfet$2_57 m1_20126_25858# vss m1_20268_25662# vss nfet$2
Xnfet$2_46 m1_20126_25858# vss m1_18073_21786# vss nfet$2
Xnfet$2_35 m1_15598_25662# m1_15822_23922# m1_16086_24542# vss nfet$2
Xnfet$2_24 m1_7095_25858# m1_7719_25662# m1_7456_23922# vss nfet$2
Xnfet$2_13 m1_11415_25662# m1_11639_23922# m1_11903_24542# vss nfet$2
Xpfet$3_7 vdd m1_354_22513# m1_354_22513# m1_n674_22102# m1_1120_21786# m1_1120_21786#
+ pfet$3
Xpfet$1_4 vdd vdd m1_3893_24224# m1_3273_23922# pfet$1
Xnfet$28_5 m1_6107_19404# m1_6107_19404# m1_n5227_21418# m1_n5227_21418# m1_n2445_21430#
+ vss nfet$28
Xpfet$1_96 vdd m1_28635_24542# vdd m1_29607_24346# pfet$1
Xpfet$1_85 vdd m1_24188_23922# m1_24452_24542# m1_23827_25858# pfet$1
Xpfet$1_74 vdd vdd m1_14556_21786# m1_15943_25858# pfet$1
Xpfet$1_63 vdd vdd m1_19781_25662# m1_19644_25858# pfet$1
Xpfet$1_52 vdd m1_20268_25662# m1_20005_23922# m1_19781_25662# pfet$1
Xpfet$1_41 vdd vdd m1_9288_21786# pd4 pfet$1
Xpfet$1_30 vdd vdd m1_2912_25858# m1_488_21786# pfet$1
Xnfet$33_3 m1_n8283_19850# m1_n8283_20611# vss vss nfet$33
Xpfet$27_4 vdd vdd m1_n5571_25662# m1_n10452_25858# pfet$27
Xnfet$6_7 m1_4005_21786# vss m1_4637_21786# vss nfet$6
Xpfet$18_0 vdd m1_32818_20470# m1_32818_20470# m1_33050_19550# m1_30256_19792# m1_30256_19792#
+ pfet$18
Xnfet$4_4 m1_9418_19550# m1_9418_19550# vss vss m1_9856_20470# vss nfet$4
Xnfet$31_0 m1_n10933_25858# m1_n8848_25658# m1_n8055_24542# vss nfet$31
Xpfet$25_1 vdd m1_n8625_26174# vdd m1_n8848_25658# pfet$25
Xnfet$5_79 m1_15921_16080# vss m1_15564_15778# vss nfet$5
Xnfet$5_68 m1_18665_17343# m1_18926_16202# m1_18441_17518# vss nfet$5
Xnfet$5_57 m1_22848_17343# m1_24904_15778# m1_24287_16080# vss nfet$5
Xnfet$5_46 m1_22034_17714# vss m1_21564_17714# vss nfet$5
Xnfet$5_24 m1_4832_17714# vss m1_1933_17343# vss nfet$5
Xnfet$5_13 m1_10458_17836# m1_11381_15778# m1_10560_16202# vss nfet$5
Xnfet$5_35 m1_n7513_20152# vss m1_5761_16080# vss nfet$5
Xnfet$10_5 m1_n789_25858# vss m1_488_21786# vss nfet$10
Xnfet$2_1 m1_2912_25858# m1_4997_25658# m1_5790_24542# vss nfet$2
Xpfet$1_109 vdd m1_12259_24224# m1_13363_25658# m1_11278_25858# pfet$1
Xnfet$2_69 m1_24309_25858# vss m1_26705_24542# vss nfet$2
Xnfet$2_58 m1_20005_23922# vss m1_20625_24224# vss nfet$2
Xnfet$2_47 m1_23964_25662# m1_24188_23922# m1_24452_24542# vss nfet$2
Xnfet$2_36 m1_11760_25858# vss m1_11039_21786# vss nfet$2
Xnfet$2_25 m1_7232_25662# m1_8076_24224# m1_9180_25658# vss nfet$2
Xnfet$2_14 m1_n7513_20152# vss m1_8692_24346# vss nfet$2
Xpfet$3_8 vdd vdd vdd m1_6360_22102# m1_5901_21590# m1_5901_21590# pfet$3
Xpfet$4_30 vdd vdd vdd m1_24560_19550# m1_21880_15478# m1_21880_15478# pfet$4
Xpfet$1_5 vdd m1_3893_24224# m1_4997_25658# m1_2912_25858# pfet$1
Xnfet$28_6 m1_n5764_21786# m1_n5764_21786# vss vss m1_n6282_21430# vss nfet$28
Xpfet$1_97 vdd vdd m1_21590_21786# m1_24309_25858# pfet$1
Xpfet$1_86 vdd m1_28634_25662# m1_28371_23922# m1_28147_25662# pfet$1
Xpfet$1_75 vdd vdd m1_19644_25858# m1_14556_21786# pfet$1
Xpfet$1_64 vdd vdd m1_22522_24542# m1_20126_25858# pfet$1
Xpfet$1_53 vdd m1_20625_24224# m1_21729_25658# m1_19644_25858# pfet$1
Xpfet$1_42 vdd m1_11760_25858# vdd m1_13363_25658# pfet$1
Xpfet$1_31 vdd m1_3273_23922# m1_3537_24542# m1_2912_25858# pfet$1
Xpfet$1_20 vdd vdd m1_4509_24346# m1_n7513_20152# pfet$1
Xpfet$27_5 vdd vdd m1_n4847_25662# m1_n10452_25858# pfet$27
Xnfet$6_8 m1_2254_21786# vss m1_2384_21590# vss nfet$6
Xpfet$18_1 vdd vdd vdd m1_33050_19550# m1_31535_19792# m1_31535_19792# pfet$18
Xnfet$24_0 m1_n6274_17836# m1_n4994_16080# m1_n5461_18030# vss nfet$24
Xnfet$31_1 m1_n10796_25662# m1_n10572_23922# m1_n10308_24542# vss nfet$31
Xpfet$25_2 vdd m1_n3651_26174# vdd m1_n4978_24224# pfet$25
.ends

.subckt nfet$47 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$45 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$44 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$42 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$40 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$48 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$46 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$44 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$43 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$41 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt asc_hysteresis_buffer$11 vss in vdd out
Xnfet$47_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$47
Xnfet$45_0 m1_348_648# vss m1_884_42# vss nfet$45
Xpfet$44_0 vdd vdd m1_884_42# m1_1156_42# pfet$44
Xpfet$42_0 vdd vdd m1_348_648# in pfet$42
Xpfet$40_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd m1_884_42#
+ m1_884_42# pfet$40
Xnfet$48_0 m1_1156_42# vss m1_884_42# vss nfet$48
Xnfet$46_0 in vss m1_348_648# vss nfet$46
Xnfet$44_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$44
Xpfet$43_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$43
Xpfet$41_0 vdd vdd m1_884_42# m1_348_648# pfet$41
.ends

.subckt pfet$69 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$67 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$73 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt nfet$71 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$70 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$68 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$74 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$72 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt asc_drive_buffer$5 vss in vdd out
Xpfet$69_0 vdd vdd m1_4002_n1060# m1_3466_n454# pfet$69
Xpfet$67_0 out out m1_4274_n1060# vdd m1_4274_n1060# out vdd vdd m1_4274_n1060# out
+ m1_4274_n1060# m1_4274_n1060# out m1_4274_n1060# vdd m1_4274_n1060# vdd m1_4274_n1060#
+ pfet$67
Xnfet$73_0 m1_3466_n454# vss m1_4002_n1060# vss nfet$73
Xnfet$71_0 m1_4274_n1060# vss m1_4002_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ m1_4274_n1060# vss m1_4002_n1060# vss nfet$71
Xpfet$70_0 vdd vdd m1_3466_n454# in pfet$70
Xpfet$68_0 m1_4274_n1060# vdd vdd m1_4274_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ vdd m1_4002_n1060# m1_4002_n1060# pfet$68
Xnfet$74_0 in vss m1_3466_n454# vss nfet$74
Xnfet$72_0 out out vss m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# m1_4274_n1060#
+ m1_4274_n1060# out m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# vss vss
+ nfet$72
.ends

.subckt xp_3_1_MUX$6 S0 S1 VDD VSS OUT_1 C_1 B_1 A_1
Xpfet$60_0 VDD A_1 m1_239_n318# m1_n432_458# pfet$60
Xpfet$60_1 VDD C_1 OUT_1 S1 pfet$60
Xpfet$60_2 VDD B_1 m1_239_n318# S0 pfet$60
Xpfet$60_3 VDD m1_239_n318# OUT_1 m1_n432_n1290# pfet$60
Xnfet$64_0 m1_n432_n1290# C_1 OUT_1 VSS nfet$64
Xnfet$64_1 m1_n432_458# B_1 m1_239_n318# VSS nfet$64
Xnfet$64_2 S1 m1_239_n318# OUT_1 VSS nfet$64
Xnfet$64_3 S0 A_1 m1_239_n318# VSS nfet$64
Xpfet$61_0 VDD VDD m1_n432_n1290# S1 pfet$61
Xpfet$61_1 VDD VDD m1_n432_458# S0 pfet$61
Xnfet$65_1 S0 VSS m1_n432_458# VSS nfet$65
Xnfet$65_0 S1 VSS m1_n432_n1290# VSS nfet$65
.ends

.subckt asc_dual_psd_def_20250809$6 vdd vss pd1 pd2 pd3 pd4 pd5 pd6 pd7 pd8 pd9 fout
+ sd1 sd2 sd3 sd4 sd5 sd6 sd7 sd8 sd9 fin define
Xnfet$4_5 m1_649_17714# m1_649_17714# vss vss m1_6971_20470# vss nfet$4
Xnfet$5_69 m1_17851_17714# vss m1_17381_17714# vss nfet$5
Xnfet$5_58 m1_23007_17836# m1_23930_15778# m1_23109_16202# vss nfet$5
Xnfet$5_47 m1_22034_17714# vss m1_22624_17518# vss nfet$5
Xnfet$10_6 m1_n910_23922# vss m1_n290_24224# vss nfet$10
Xnfet$5_25 m1_2092_17836# m1_3372_16080# m1_2905_18030# vss nfet$5
Xnfet$5_14 m1_6116_17343# m1_8172_15778# m1_7555_16080# vss nfet$5
Xnfet$5_36 m1_n3064_17714# vss m1_n2474_17518# vss nfet$5
Xpfet$30_0 vdd m1_n6380_21786# m1_n6380_21786# m1_n5019_19550# m1_n5227_20152# m1_n5227_20152#
+ pfet$30
Xnfet$2_2 m1_n7513_20152# vss m1_4509_24346# vss nfet$2
Xnfet$2_59 m1_19644_25858# m1_20268_25662# m1_20005_23922# vss nfet$2
Xnfet$2_48 m1_18073_21786# vss m1_23827_25858# vss nfet$2
Xnfet$2_37 m1_11039_21786# vss m1_15461_25858# vss nfet$2
Xnfet$2_26 m1_7095_25858# m1_9180_25658# m1_9973_24542# vss nfet$2
Xnfet$2_15 m1_7232_25662# m1_7456_23922# m1_7720_24542# vss nfet$2
Xpfet$4_31 vdd m1_n2543_20130# m1_n2543_20130# m1_20407_19850# m1_19969_19550# m1_19969_19550#
+ pfet$4
Xpfet$4_20 vdd m1_n3822_21786# m1_n3822_21786# m1_14009_19550# m1_9015_17714# m1_9015_17714#
+ pfet$4
Xpfet$3_9 vdd m1_3871_22513# m1_3871_22513# m1_3471_22402# m1_4005_21786# m1_4005_21786#
+ pfet$3
Xpfet$1_6 vdd vdd m1_3536_25662# m1_3394_25858# pfet$1
Xnfet$28_7 m1_n3822_21786# m1_n3822_21786# m1_n4485_21904# m1_n4485_21904# m1_n3724_21430#
+ vss nfet$28
Xpfet$1_65 vdd vdd m1_18073_21786# m1_20126_25858# pfet$1
Xpfet$1_54 vdd vdd m1_24808_24224# m1_24188_23922# pfet$1
Xpfet$1_43 vdd vdd m1_12805_21786# pd5 pfet$1
Xpfet$1_32 vdd vdd m1_7720_24542# m1_8076_24224# pfet$1
Xpfet$1_21 vdd m1_7456_23922# m1_7720_24542# m1_7095_25858# pfet$1
Xpfet$1_10 vdd m1_8076_24224# m1_9180_25658# m1_7095_25858# pfet$1
Xpfet$27_6 vdd vdd m1_n4623_25487# fin pfet$27
Xpfet$1_98 vdd m1_30095_25658# m1_30888_24542# m1_28147_25662# pfet$1
Xpfet$1_87 vdd vdd m1_28147_25662# m1_28010_25858# pfet$1
Xpfet$1_76 vdd m1_20005_23922# m1_20269_24542# m1_19644_25858# pfet$1
Xnfet$6_9 m1_23356_21786# vss m1_23486_21590# vss nfet$6
Xpfet$18_2 vdd m1_32818_21586# m1_32818_21586# m1_33050_22344# m1_30256_22102# m1_30256_22102#
+ pfet$18
Xnfet$17_0 m1_31535_22102# m1_32818_21586# vss vss nfet$17
Xnfet$24_1 m1_n6433_17343# m1_n4377_15778# m1_n4994_16080# vss nfet$24
Xnfet$31_2 m1_n10933_25858# m1_n10309_25662# m1_n10572_23922# vss nfet$31
Xpfet$25_3 vdd vdd m1_n3651_26174# m1_n3541_23922# pfet$25
Xnfet$4_6 m1_n1133_19550# m1_n1133_19550# vss vss m1_n695_20470# vss nfet$4
Xnfet$10_7 m1_25107_21786# vss m1_32193_25858# vss nfet$10
Xnfet$5_59 m1_17851_17714# vss m1_20721_15778# vss nfet$5
Xnfet$5_48 m1_18824_17836# m1_20104_16080# m1_19637_18030# vss nfet$5
Xnfet$5_26 m1_5302_17714# vss m1_5892_17518# vss nfet$5
Xnfet$5_15 m1_5302_17714# vss m1_8172_15778# vss nfet$5
Xnfet$5_37 m1_n7513_20152# vss m1_n2605_16080# vss nfet$5
Xpfet$30_1 vdd vdd vdd m1_n5019_22344# m1_n4485_21904# m1_n4485_21904# pfet$30
Xpfet$23_0 vdd m1_n10309_25662# m1_n10572_23922# m1_n10796_25662# pfet$23
Xnfet$2_3 m1_488_21786# vss m1_2912_25858# vss nfet$2
Xnfet$2_49 m1_19781_25662# m1_20005_23922# m1_20269_24542# vss nfet$2
Xnfet$2_38 m1_n7513_20152# vss m1_12875_24346# vss nfet$2
Xnfet$2_27 m1_7577_25858# vss m1_7719_25662# vss nfet$2
Xnfet$2_16 m1_4005_21786# vss m1_7095_25858# vss nfet$2
Xpfet$4_32 vdd m1_n2543_20130# m1_n2543_20130# m1_21043_19550# m1_17381_17714# m1_17381_17714#
+ pfet$4
Xpfet$4_21 vdd vdd vdd m1_13373_19850# m1_15171_20152# m1_15171_20152# pfet$4
Xpfet$4_10 vdd vdd vdd m1_9856_19850# m1_11654_20152# m1_11654_20152# pfet$4
Xpfet$8_0 vdd vdd m1_n7401_15478# sd9 pfet$8
Xnfet$28_8 m1_9624_19404# m1_9624_19404# vss vss m1_n3724_21430# vss nfet$28
Xpfet$1_7 vdd vdd m1_7232_25662# m1_7095_25858# pfet$1
Xpfet$1_99 vdd vdd m1_26705_24542# m1_24309_25858# pfet$1
Xpfet$1_88 vdd vdd m1_28634_25662# m1_28492_25858# pfet$1
Xpfet$1_77 vdd vdd m1_20269_24542# m1_20625_24224# pfet$1
Xpfet$1_66 vdd vdd m1_15461_25858# m1_11039_21786# pfet$1
Xpfet$1_55 vdd m1_24451_25662# m1_24188_23922# m1_23964_25662# pfet$1
Xpfet$1_44 vdd m1_15943_25858# vdd m1_17546_25658# pfet$1
Xpfet$1_33 vdd vdd m1_7522_21786# m1_7577_25858# pfet$1
Xpfet$1_22 vdd vdd m1_3537_24542# m1_3893_24224# pfet$1
Xpfet$1_11 vdd vdd m1_7719_25662# m1_7577_25858# pfet$1
Xpfet$27_7 vdd vdd m1_n3541_23922# m1_n3184_24224# pfet$27
Xnfet$24_2 m1_n6274_17836# m1_n5351_15778# m1_n6172_16202# vss nfet$24
Xnfet$31_3 m1_n10796_25662# m1_n9952_24224# m1_n8848_25658# vss nfet$31
Xpfet$25_4 vdd m1_n10452_25858# vdd m1_n4362_24346# pfet$25
Xnfet$4_7 m1_n7383_17599# m1_n7383_17599# vss vss m1_n63_20470# vss nfet$4
Xnfet$10_8 m1_32193_25858# vss m1_32330_25662# vss nfet$10
Xnfet$5_49 m1_21564_17714# vss m1_18665_17343# vss nfet$5
Xpfet$7_10 vdd vdd m1_29239_20152# m1_26063_15478# pfet$7
Xnfet$5_27 m1_1119_17714# vss m1_3989_15778# vss nfet$5
Xnfet$5_16 m1_6275_17836# m1_7198_15778# m1_6377_16202# vss nfet$5
Xnfet$5_38 m1_n2250_17343# m1_n1989_16202# m1_n2474_17518# vss nfet$5
Xpfet$16_0 vdd vdd vdd m1_36073_22344# define define pfet$16
Xpfet$30_2 vdd m1_n5764_21786# m1_n5764_21786# m1_n5019_22344# m1_n5227_21418# m1_n5227_21418#
+ pfet$30
Xpfet$23_1 vdd m1_n9952_24224# m1_n8848_25658# m1_n10933_25858# pfet$23
Xnfet$2_4 m1_2912_25858# vss m1_3049_25662# vss nfet$2
Xnfet$29_10 vss vss m1_n4978_24224# vss nfet$29
Xnfet$2_39 pd4 vss m1_9288_21786# vss nfet$2
Xpfet$4_33 vdd m1_n3206_20274# m1_n3206_20274# m1_24560_19550# m1_21564_17714# m1_21564_17714#
+ pfet$4
Xpfet$4_22 vdd vdd vdd m1_14009_19550# m1_9331_15478# m1_9331_15478# pfet$4
Xnfet$2_28 m1_3394_25858# vss m1_4005_21786# vss nfet$2
Xnfet$2_17 m1_11639_23922# vss m1_12259_24224# vss nfet$2
Xpfet$4_11 vdd vdd vdd m1_10492_19550# m1_5148_15478# m1_5148_15478# pfet$4
Xpfet$8_1 vdd vdd m1_21880_15478# sd2 pfet$8
Xnfet$28_9 m1_n6380_21786# m1_n6380_21786# m1_n6839_21786# m1_n6839_21786# m1_n6282_21430#
+ vss nfet$28
Xpfet$1_8 vdd vdd m1_8076_24224# m1_7456_23922# pfet$1
Xpfet$1_89 vdd vdd m1_19839_21786# pd7 pfet$1
Xpfet$1_78 vdd m1_20269_24542# vdd m1_21241_24346# pfet$1
Xpfet$1_67 vdd m1_15822_23922# m1_16086_24542# m1_15461_25858# pfet$1
Xpfet$1_56 vdd m1_24808_24224# m1_25912_25658# m1_23827_25858# pfet$1
Xpfet$1_45 vdd vdd m1_16442_24224# m1_15822_23922# pfet$1
Xpfet$1_34 vdd m1_9180_25658# m1_9973_24542# m1_7232_25662# pfet$1
Xpfet$1_23 vdd m1_3537_24542# vdd m1_4509_24346# pfet$1
Xpfet$1_12 vdd m1_7577_25858# vdd m1_9180_25658# pfet$1
Xpfet$27_8 vdd vdd m1_n2567_23922# m1_n7320_25516# pfet$27
Xpfet$25_5 vdd vdd m1_n10308_24542# m1_n9952_24224# pfet$25
Xnfet$4_8 m1_27003_19550# m1_27003_19550# vss vss m1_27441_20470# vss nfet$4
Xnfet$24_3 m1_n6433_17343# m1_n6172_16202# m1_n6657_17518# vss nfet$24
Xnfet$31_4 m1_n4623_25487# m1_n2567_23922# m1_n3184_24224# vss nfet$31
Xnfet$10_9 m1_n7513_20152# vss m1_33790_24346# vss nfet$10
Xnfet$5_28 m1_1933_17343# vss m1_2092_17836# vss nfet$5
Xnfet$5_17 m1_649_17714# vss m1_n2250_17343# vss nfet$5
Xnfet$5_39 m1_n3064_17714# vss m1_n3534_17714# vss nfet$5
Xpfet$16_1 vdd m1_35837_22102# m1_35837_22102# m1_36073_22344# fout fout pfet$16
Xpfet$7_11 vdd vdd m1_18688_20152# m1_13514_15478# pfet$7
Xnfet$22_0 m1_4620_20152# m1_4620_20152# m1_2590_19404# m1_2590_19404# m1_3454_20470#
+ vss nfet$22
Xpfet$23_2 vdd m1_n4362_24346# m1_n4847_25662# m1_n4464_25980# pfet$23
Xnfet$2_5 m1_2912_25858# m1_3536_25662# m1_3273_23922# vss nfet$2
Xnfet$29_11 m1_n10452_25858# vss m1_n4847_25662# vss nfet$29
Xnfet$2_29 m1_15943_25858# vss m1_14556_21786# vss nfet$2
Xpfet$4_34 vdd m1_n3206_20274# m1_n3206_20274# m1_23924_19850# m1_23486_19550# m1_23486_19550#
+ pfet$4
Xpfet$4_23 vdd vdd vdd m1_16890_19850# m1_18688_20152# m1_18688_20152# pfet$4
Xnfet$2_18 m1_7095_25858# vss m1_7232_25662# vss nfet$2
Xpfet$4_12 vdd m1_6107_19404# m1_6107_19404# m1_6975_19550# m1_649_17714# m1_649_17714#
+ pfet$4
Xpfet$8_2 vdd vdd m1_26063_15478# sd1 pfet$8
Xpfet$1_9 vdd m1_7719_25662# m1_7456_23922# m1_7232_25662# pfet$1
Xpfet$1_79 vdd m1_17546_25658# m1_18339_24542# m1_15598_25662# pfet$1
Xpfet$1_68 vdd vdd m1_16086_24542# m1_16442_24224# pfet$1
Xpfet$1_57 vdd vdd m1_24451_25662# m1_24309_25858# pfet$1
Xpfet$1_46 vdd m1_16442_24224# m1_17546_25658# m1_15461_25858# pfet$1
Xpfet$1_35 vdd m1_7720_24542# vdd m1_8692_24346# pfet$1
Xpfet$1_24 vdd vdd m1_5790_24542# m1_3394_25858# pfet$1
Xpfet$1_13 vdd vdd m1_12259_24224# m1_11639_23922# pfet$1
Xpfet$27_9 vdd vdd m1_n4464_25980# m1_n4623_25487# pfet$27
Xnfet$4_9 m1_25747_17714# m1_25747_17714# vss vss m1_28073_20470# vss nfet$4
Xnfet$24_4 m1_27031_17343# m1_27292_16202# m1_26807_17518# vss nfet$24
Xnfet$31_5 m1_n4464_25980# m1_n3541_23922# m1_n4362_24346# vss nfet$31
Xpfet$25_6 vdd m1_n10308_24542# vdd m1_n9336_24346# pfet$25
Xnfet$5_29 m1_3372_16080# vss m1_3015_15778# vss nfet$5
Xnfet$5_18 m1_1119_17714# vss m1_649_17714# vss nfet$5
Xpfet$7_12 vdd vdd m1_15171_20152# m1_9331_15478# pfet$7
Xnfet$22_1 m1_1103_20152# m1_1103_20152# m1_n927_19404# m1_n927_19404# m1_n63_20470#
+ vss nfet$22
Xpfet$23_3 vdd m1_n3184_24224# m1_n3651_26174# m1_n4623_25487# pfet$23
Xnfet$15_0 m1_21456_22513# m1_21456_22513# m1_30256_19792# m1_30256_19792# m1_30492_20470#
+ vss nfet$15
Xnfet$2_6 m1_3049_25662# m1_3893_24224# m1_4997_25658# vss nfet$2
Xnfet$29_12 m1_n10452_25858# vss m1_n5571_25662# vss nfet$29
Xpfet$21_0 vdd vdd m1_n7513_20152# m1_35837_22102# pfet$21
Xnfet$2_19 m1_7456_23922# vss m1_8076_24224# vss nfet$2
Xpfet$4_35 vdd m1_n3822_21786# m1_n3822_21786# m1_13373_19850# m1_12935_19550# m1_12935_19550#
+ pfet$4
Xpfet$4_24 vdd m1_n1927_20274# m1_n1927_20274# m1_16890_19850# m1_16452_19550# m1_16452_19550#
+ pfet$4
Xpfet$4_13 vdd m1_n927_19404# m1_n927_19404# m1_n695_19850# m1_n1133_19550# m1_n1133_19550#
+ pfet$4
Xpfet$6_0 vdd vdd m1_n6274_17836# m1_n6433_17343# pfet$6
Xpfet$1_69 vdd vdd m1_12875_24346# m1_n7513_20152# pfet$1
Xpfet$1_58 vdd vdd m1_23964_25662# m1_23827_25858# pfet$1
Xpfet$1_47 vdd vdd m1_15943_25858# m1_17058_24346# pfet$1
Xpfet$1_36 vdd vdd m1_8692_24346# m1_n7513_20152# pfet$1
Xpfet$1_25 vdd vdd m1_4005_21786# m1_3394_25858# pfet$1
Xpfet$1_14 vdd vdd m1_11902_25662# m1_11760_25858# pfet$1
Xnfet$24_5 m1_27031_17343# m1_29087_15778# m1_28470_16080# vss nfet$24
Xnfet$31_6 m1_n4464_25980# m1_n3184_24224# m1_n3651_26174# vss nfet$31
Xpfet$25_7 vdd vdd m1_n10452_25858# m1_n4978_24224# pfet$25
Xpfet$2_90 vdd m1_19747_15778# m1_18926_16202# m1_18665_17343# pfet$2
Xnfet$9_0 m1_n3534_17714# vss m1_n6433_17343# vss nfet$9
Xpfet$7_13 vdd vdd m1_16452_19550# m1_13198_17714# pfet$7
Xnfet$5_19 m1_n7513_20152# vss m1_1578_16080# vss nfet$5
Xpfet$23_4 vdd m1_n2567_23922# m1_n3184_24224# m1_n4464_25980# pfet$23
Xnfet$15_1 m1_14422_22513# m1_14422_22513# m1_31535_19792# m1_31535_19792# m1_31771_20470#
+ vss nfet$15
Xnfet$2_7 m1_3049_25662# m1_3273_23922# m1_3537_24542# vss nfet$2
Xnfet$22_2 m1_n3218_15478# m1_n3218_15478# m1_2590_19404# m1_2590_19404# m1_2822_20470#
+ vss nfet$22
Xnfet$29_13 fin vss m1_n4623_25487# vss nfet$29
Xpfet$14_0 vdd vdd m1_n1263_21786# pd1 pfet$14
Xpfet$4_25 vdd vdd vdd m1_17526_19550# m1_13514_15478# m1_13514_15478# pfet$4
Xpfet$4_14 vdd m1_n927_19404# m1_n927_19404# m1_n59_19550# m1_n7383_17599# m1_n7383_17599#
+ pfet$4
Xpfet$6_1 vdd vdd m1_n4377_15778# m1_n7247_17714# pfet$6
Xpfet$1_59 vdd vdd m1_16322_21786# pd6 pfet$1
Xpfet$1_48 vdd m1_16085_25662# m1_15822_23922# m1_15598_25662# pfet$1
Xpfet$1_37 vdd vdd m1_9973_24542# m1_7577_25858# pfet$1
Xpfet$1_26 vdd m1_4997_25658# m1_5790_24542# m1_3049_25662# pfet$1
Xpfet$1_15 vdd m1_11902_25662# m1_11639_23922# m1_11415_25662# pfet$1
Xnfet$24_6 m1_27190_17836# m1_28113_15778# m1_27292_16202# vss nfet$24
Xnfet$31_7 m1_n4623_25487# m1_n4362_24346# m1_n4847_25662# vss nfet$31
Xpfet$2_91 vdd m1_24287_16080# m1_23820_18030# m1_22848_17343# pfet$2
Xpfet$2_80 vdd vdd m1_15564_15778# m1_15921_16080# pfet$2
Xpfet$7_14 vdd vdd m1_23486_19550# m1_21564_17714# pfet$7
Xnfet$9_1 m1_n7513_20152# vss m1_n6788_16080# vss nfet$9
Xnfet$15_2 m1_17939_22513# m1_17939_22513# vss vss m1_31771_20470# vss nfet$15
Xnfet$2_8 m1_3394_25858# vss m1_3536_25662# vss nfet$2
Xnfet$22_3 m1_8137_20152# m1_8137_20152# m1_6107_19404# m1_6107_19404# m1_6971_20470#
+ vss nfet$22
Xpfet$23_5 vdd m1_n10572_23922# m1_n10308_24542# m1_n10933_25858# pfet$23
Xpfet$14_1 vdd vdd m1_2254_21786# pd2 pfet$14
Xnfet$20_0 fout vss m1_35837_22102# vss nfet$20
Xpfet$4_26 vdd m1_n1927_20274# m1_n1927_20274# m1_17526_19550# m1_13198_17714# m1_13198_17714#
+ pfet$4
Xpfet$4_15 vdd vdd vdd m1_n59_19550# m1_n7401_15478# m1_n7401_15478# pfet$4
Xpfet$6_2 vdd vdd m1_n5351_15778# m1_n4994_16080# pfet$6
Xpfet$1_49 vdd m1_20126_25858# vdd m1_21729_25658# pfet$1
Xpfet$1_38 vdd vdd m1_16085_25662# m1_15943_25858# pfet$1
Xpfet$1_27 vdd vdd m1_11278_25858# m1_7522_21786# pfet$1
Xpfet$1_16 vdd vdd m1_5771_21786# pd3 pfet$1
Xnfet$24_7 m1_27190_17836# m1_28470_16080# m1_28003_18030# vss nfet$24
Xpfet$2_92 vdd m1_15454_18030# vdd m1_14127_16080# pfet$2
Xpfet$2_81 vdd vdd m1_13668_17714# m1_14127_16080# pfet$2
Xpfet$2_70 vdd vdd m1_18824_17836# m1_18665_17343# pfet$2
Xpfet$7_15 vdd vdd m1_22205_20152# m1_17697_15478# pfet$7
Xnfet$9_2 m1_n4994_16080# vss m1_n5351_15778# vss nfet$9
Xnfet$15_3 m1_24973_22513# m1_24973_22513# vss vss m1_30492_20470# vss nfet$15
Xnfet$22_4 m1_965_15478# m1_965_15478# m1_6107_19404# m1_6107_19404# m1_6339_20470#
+ vss nfet$22
Xpfet$23_6 vdd m1_n8848_25658# m1_n8055_24542# m1_n10796_25662# pfet$23
Xnfet$2_9 m1_3273_23922# vss m1_3893_24224# vss nfet$2
Xpfet$14_2 vdd vdd m1_26873_21786# pd9 pfet$14
Xnfet$20_1 define m1_35837_22102# vss vss nfet$20
Xnfet$13_0 m1_n290_24224# m1_n290_24224# m1_n646_24542# m1_n646_24542# m1_n192_24542#
+ vss nfet$13
Xpfet$4_27 vdd vdd vdd m1_20407_19850# m1_22205_20152# m1_22205_20152# pfet$4
Xpfet$4_16 vdd vdd vdd m1_28077_19550# m1_26063_15478# m1_26063_15478# pfet$4
Xnfet$3_10 m1_19839_21786# m1_19839_21786# m1_21456_22513# m1_21456_22513# m1_21060_21586#
+ vss nfet$3
Xpfet$6_3 vdd vdd m1_n6657_17518# m1_n7247_17714# pfet$6
Xpfet$1_39 vdd vdd m1_15598_25662# m1_15461_25858# pfet$1
Xpfet$1_28 vdd m1_11639_23922# m1_11903_24542# m1_11278_25858# pfet$1
Xpfet$1_17 vdd vdd m1_7577_25858# m1_8692_24346# pfet$1
Xpfet$4_0 vdd m1_2590_19404# m1_2590_19404# m1_3458_19550# m1_n3534_17714# m1_n3534_17714#
+ pfet$4
Xpfet$2_93 vdd m1_23820_18030# vdd m1_22493_16080# pfet$2
Xpfet$2_82 vdd m1_13668_17714# vdd m1_14743_16202# pfet$2
Xpfet$2_71 vdd vdd m1_19747_15778# m1_20104_16080# pfet$2
Xpfet$2_60 vdd vdd m1_n194_15778# m1_n3064_17714# pfet$2
Xnfet$9_3 m1_n6433_17343# vss m1_n6274_17836# vss nfet$9
Xpfet$7_16 vdd vdd m1_19969_19550# m1_17381_17714# pfet$7
Xnfet$15_4 m1_32818_20470# m1_32818_20470# vss vss m1_34329_20470# vss nfet$15
Xnfet$22_5 m1_5148_15478# m1_5148_15478# m1_9624_19404# m1_9624_19404# m1_9856_20470#
+ vss nfet$22
Xpfet$23_7 vdd m1_n3541_23922# m1_n4362_24346# m1_n4623_25487# pfet$23
Xnfet$7_0 m1_n3534_17714# vss m1_2384_19550# vss nfet$7
Xnfet$6_10 m1_21590_21786# vss m1_22222_21786# vss nfet$6
Xnfet$13_1 m1_814_25658# m1_814_25658# vss vss m1_1273_25502# vss nfet$13
Xpfet$4_28 vdd vdd vdd m1_21043_19550# m1_17697_15478# m1_17697_15478# pfet$4
Xpfet$4_17 vdd m1_n3822_20130# m1_n3822_20130# m1_28077_19550# m1_25747_17714# m1_25747_17714#
+ pfet$4
Xpfet$12_0 vdd m1_31535_19792# vdd m1_17939_22513# pfet$12
Xnfet$3_11 m1_19969_21590# m1_19969_21590# m1_21456_22513# m1_21456_22513# m1_20428_21586#
+ vss nfet$3
Xpfet$6_4 vdd vdd m1_n6433_17343# m1_n3534_17714# pfet$6
Xpfet$1_29 vdd vdd m1_11903_24542# m1_12259_24224# pfet$1
Xpfet$1_18 vdd vdd m1_11415_25662# m1_11278_25858# pfet$1
Xpfet$4_1 vdd vdd vdd m1_2822_19850# m1_4620_20152# m1_4620_20152# pfet$4
Xnfet$9_10 m1_26217_17714# vss m1_29087_15778# vss nfet$9
Xpfet$2_94 vdd vdd m1_22624_17518# m1_22034_17714# pfet$2
Xpfet$2_83 vdd m1_16538_15778# m1_15921_16080# m1_14641_17836# pfet$2
Xpfet$2_72 vdd m1_20721_15778# m1_20104_16080# m1_18824_17836# pfet$2
Xpfet$2_61 vdd m1_n811_16080# m1_n1278_18030# m1_n2250_17343# pfet$2
Xpfet$2_50 vdd m1_n1168_15778# m1_n1989_16202# m1_n2250_17343# pfet$2
Xnfet$9_4 m1_n7247_17714# vss m1_n4377_15778# vss nfet$9
Xnfet$36_0 m1_n4485_20152# m1_n6380_21786# vss vss nfet$36
Xpfet$7_17 vdd vdd m1_25722_20152# m1_21880_15478# pfet$7
Xnfet$22_6 m1_11654_20152# m1_11654_20152# m1_9624_19404# m1_9624_19404# m1_10488_20470#
+ vss nfet$22
Xnfet$15_5 m1_32818_21586# m1_32818_21586# m1_34093_19792# m1_34093_19792# m1_34329_20470#
+ vss nfet$15
Xnfet$7_1 m1_n3218_15478# vss m1_4620_20152# vss nfet$7
Xnfet$6_11 m1_18073_21786# vss m1_18705_21786# vss nfet$6
Xnfet$13_2 m1_326_24346# m1_326_24346# m1_n789_25858# m1_n789_25858# m1_1273_25502#
+ vss nfet$13
Xpfet$4_29 vdd vdd vdd m1_23924_19850# m1_25722_20152# m1_25722_20152# pfet$4
Xpfet$4_18 vdd vdd vdd m1_27441_19850# m1_29239_20152# m1_29239_20152# pfet$4
Xpfet$12_1 vdd vdd m1_30256_19792# m1_21456_22513# pfet$12
Xnfet$3_12 m1_16322_21786# m1_16322_21786# m1_17939_22513# m1_17939_22513# m1_17543_21586#
+ vss nfet$3
Xpfet$6_5 vdd vdd m1_n6788_16080# m1_n7513_20152# pfet$6
Xpfet$1_19 vdd vdd m1_7095_25858# m1_4005_21786# pfet$1
Xpfet$4_2 vdd m1_2590_19404# m1_2590_19404# m1_2822_19850# m1_2384_19550# m1_2384_19550#
+ pfet$4
Xnfet$9_11 m1_27031_17343# vss m1_27190_17836# vss nfet$9
Xpfet$2_95 vdd vdd m1_21564_17714# m1_22034_17714# pfet$2
Xpfet$2_84 vdd vdd m1_17381_17714# m1_17851_17714# pfet$2
Xpfet$2_73 vdd vdd m1_16538_15778# m1_13668_17714# pfet$2
Xpfet$2_62 vdd vdd m1_23007_17836# m1_22848_17343# pfet$2
Xpfet$2_40 vdd m1_10560_16202# m1_10075_17518# m1_10458_17836# pfet$2
Xpfet$2_51 vdd vdd m1_n1168_15778# m1_n811_16080# pfet$2
Xnfet$9_5 m1_n7247_17714# vss m1_n6657_17518# vss nfet$9
Xnfet$36_1 m1_n5227_20152# vss m1_n6380_21786# vss nfet$36
Xnfet$29_0 m1_n8625_26174# vss m1_n8055_24542# vss nfet$29
Xnfet$15_6 m1_354_22513# m1_354_22513# m1_31535_22102# m1_31535_22102# m1_31771_21430#
+ vss nfet$15
Xnfet$22_7 m1_n7401_15478# m1_n7401_15478# m1_n927_19404# m1_n927_19404# m1_n695_20470#
+ vss nfet$22
Xnfet$7_2 m1_n7401_15478# vss m1_1103_20152# vss nfet$7
Xnfet$6_12 m1_14556_21786# vss m1_15188_21786# vss nfet$6
Xnfet$13_3 m1_326_24346# m1_326_24346# vss vss m1_n192_24542# vss nfet$13
Xpfet$4_19 vdd m1_n3822_20130# m1_n3822_20130# m1_27441_19850# m1_27003_19550# m1_27003_19550#
+ pfet$4
Xpfet$12_2 vdd m1_30256_19792# vdd m1_24973_22513# pfet$12
Xnfet$11_0 m1_n1134_25662# m1_n910_23922# m1_n646_24542# vss nfet$11
Xnfet$3_13 m1_16452_21590# m1_16452_21590# m1_17939_22513# m1_17939_22513# m1_16911_21586#
+ vss nfet$3
Xpfet$6_6 vdd vdd m1_n7383_17599# m1_n7247_17714# pfet$6
Xpfet$4_3 vdd vdd vdd m1_3458_19550# m1_n3218_15478# m1_n3218_15478# pfet$4
Xpfet$2_96 vdd vdd m1_18665_17343# m1_21564_17714# pfet$2
Xpfet$2_85 vdd m1_18926_16202# m1_18441_17518# m1_18824_17836# pfet$2
Xpfet$2_74 vdd vdd m1_14641_17836# m1_14482_17343# pfet$2
Xpfet$2_63 vdd m1_23930_15778# m1_23109_16202# m1_22848_17343# pfet$2
Xnfet$9_12 m1_28470_16080# vss m1_28113_15778# vss nfet$9
Xpfet$2_30 vdd vdd m1_1933_17343# m1_4832_17714# pfet$2
Xpfet$2_41 vdd vdd m1_10075_17518# m1_9485_17714# pfet$2
Xpfet$2_52 vdd m1_n3064_17714# vdd m1_n1989_16202# pfet$2
Xnfet$29_1 m1_n8625_26174# vss m1_n7082_23622# vss nfet$29
Xpfet$2_0 vdd vdd m1_12355_15778# m1_9485_17714# pfet$2
Xnfet$9_6 m1_n7247_17714# vss m1_n7383_17599# vss nfet$9
Xnfet$15_7 m1_3871_22513# m1_3871_22513# vss vss m1_31771_21430# vss nfet$15
Xnfet$22_8 m1_26063_15478# m1_26063_15478# m1_n3822_20130# m1_n3822_20130# m1_27441_20470#
+ vss nfet$22
Xnfet$10_10 m1_32675_25947# vss m1_35071_24542# vss nfet$10
Xnfet$7_3 m1_649_17714# vss m1_5901_19550# vss nfet$7
Xpfet$28_0 vdd vdd m1_n7186_25858# m1_n10452_25858# pfet$28
Xnfet$6_13 m1_16322_21786# vss m1_16452_21590# vss nfet$6
Xnfet$13_4 m1_33174_24224# m1_33174_24224# m1_32818_24542# m1_32818_24542# m1_33272_24542#
+ vss nfet$13
Xnfet$21_20 m1_22493_16080# m1_22493_16080# m1_22034_17714# m1_22034_17714# m1_22591_16398#
+ vss nfet$21
Xnfet$5_0 m1_9485_17714# vss m1_9015_17714# vss nfet$5
Xpfet$12_3 vdd vdd m1_34843_21786# m1_34093_19792# pfet$12
Xnfet$11_1 m1_n1271_25858# m1_n647_25662# m1_n910_23922# vss nfet$11
Xnfet$3_14 m1_12805_21786# m1_12805_21786# m1_14422_22513# m1_14422_22513# m1_14026_21586#
+ vss nfet$3
Xpfet$6_7 vdd vdd m1_27190_17836# m1_27031_17343# pfet$6
Xpfet$10_0 vdd vdd m1_n646_24542# m1_n290_24224# pfet$10
Xpfet$4_4 vdd m1_6107_19404# m1_6107_19404# m1_6339_19850# m1_5901_19550# m1_5901_19550#
+ pfet$4
Xnfet$9_13 m1_26217_17714# vss m1_25747_17714# vss nfet$9
Xpfet$2_97 vdd vdd m1_22493_16080# m1_n7513_20152# pfet$2
Xpfet$2_86 vdd m1_19637_18030# vdd m1_18310_16080# pfet$2
Xpfet$2_75 vdd vdd m1_17697_15478# sd3 pfet$2
Xpfet$2_64 vdd vdd m1_23930_15778# m1_24287_16080# pfet$2
Xpfet$2_20 vdd vdd m1_1119_17714# m1_1578_16080# pfet$2
Xpfet$2_31 vdd m1_3372_16080# m1_2905_18030# m1_1933_17343# pfet$2
Xpfet$2_42 vdd m1_11271_18030# vdd m1_9944_16080# pfet$2
Xpfet$2_53 vdd vdd m1_n3218_15478# sd8 pfet$2
Xnfet$29_2 vss vss m1_n9336_24346# vss nfet$29
Xnfet$9_7 m1_26217_17714# vss m1_26807_17518# vss nfet$9
Xpfet$2_1 vdd vdd m1_11381_15778# m1_11738_16080# pfet$2
Xnfet$22_9 m1_29239_20152# m1_29239_20152# m1_n3822_20130# m1_n3822_20130# m1_28073_20470#
+ vss nfet$22
Xnfet$10_11 m1_32554_23922# vss m1_33174_24224# vss nfet$10
Xnfet$34_0 m1_n4485_21904# m1_n5764_21786# vss vss nfet$34
Xpfet$28_1 vdd m1_n7186_25858# vdd m1_n6111_25858# pfet$28
Xnfet$6_14 m1_19839_21786# vss m1_19969_21590# vss nfet$6
Xnfet$7_4 m1_4832_17714# vss m1_9418_19550# vss nfet$7
Xnfet$13_5 m1_33790_24346# m1_33790_24346# vss vss m1_33272_24542# vss nfet$13
Xnfet$21_21 m1_14127_16080# m1_14127_16080# vss vss m1_15690_17358# vss nfet$21
Xnfet$21_10 m1_1578_16080# m1_1578_16080# m1_1119_17714# m1_1119_17714# m1_1676_16398#
+ vss nfet$21
Xnfet$5_1 m1_9015_17714# vss m1_6116_17343# vss nfet$5
Xpfet$12_4 vdd m1_34093_19792# vdd m1_32818_20470# pfet$12
Xnfet$11_2 m1_n1271_25858# m1_814_25658# m1_1607_24542# vss nfet$11
Xnfet$3_15 m1_26873_21786# m1_26873_21786# m1_28490_22513# m1_28490_22513# m1_28094_21586#
+ vss nfet$3
Xpfet$6_8 vdd vdd m1_28113_15778# m1_28470_16080# pfet$6
Xpfet$10_1 vdd m1_n789_25858# vdd m1_814_25658# pfet$10
Xpfet$4_5 vdd vdd vdd m1_n695_19850# m1_1103_20152# m1_1103_20152# pfet$4
Xpfet$2_98 vdd m1_20104_16080# m1_19637_18030# m1_18665_17343# pfet$2
Xpfet$2_87 vdd vdd m1_18310_16080# m1_n7513_20152# pfet$2
Xpfet$2_76 vdd m1_17851_17714# vdd m1_18926_16202# pfet$2
Xpfet$2_65 vdd m1_24904_15778# m1_24287_16080# m1_23007_17836# pfet$2
Xpfet$2_21 vdd vdd m1_965_15478# sd7 pfet$2
Xpfet$2_10 vdd m1_8172_15778# m1_7555_16080# m1_6275_17836# pfet$2
Xpfet$2_32 vdd vdd m1_2905_18030# m1_3015_15778# pfet$2
Xpfet$2_43 vdd vdd m1_11271_18030# m1_11381_15778# pfet$2
Xpfet$2_54 vdd vdd m1_n1278_18030# m1_n1168_15778# pfet$2
Xnfet$29_3 fin vss m1_n10933_25858# vss nfet$29
Xnfet$9_8 m1_n7513_20152# vss m1_26676_16080# vss nfet$9
Xpfet$2_2 vdd m1_12355_15778# m1_11738_16080# m1_10458_17836# pfet$2
Xnfet$10_12 m1_32675_25947# vss m1_28624_21786# vss nfet$10
Xnfet$34_1 m1_n5227_21418# vss m1_n5764_21786# vss nfet$34
Xnfet$27_0 m1_n7082_23622# m1_n6856_24542# vss vss nfet$27
Xnfet$7_5 m1_965_15478# vss m1_8137_20152# vss nfet$7
Xnfet$13_6 m1_33790_24346# m1_33790_24346# m1_32675_25947# m1_32675_25947# m1_34737_25502#
+ vss nfet$13
Xnfet$6_15 m1_28624_21786# vss m1_29256_21786# vss nfet$6
Xnfet$21_22 m1_15564_15778# m1_15564_15778# m1_15454_18030# m1_15454_18030# m1_15690_17358#
+ vss nfet$21
Xnfet$5_2 m1_6275_17836# m1_7555_16080# m1_7088_18030# vss nfet$5
Xnfet$21_11 m1_6377_16202# m1_6377_16202# vss vss m1_5859_16398# vss nfet$21
Xpfet$33_0 vdd vdd m1_n8145_21908# m1_n6839_20152# pfet$33
Xpfet$12_5 vdd vdd m1_34093_19792# m1_32818_21586# pfet$12
Xnfet$11_3 m1_n1134_25662# m1_n290_24224# m1_814_25658# vss nfet$11
Xnfet$3_16 m1_27003_21590# m1_27003_21590# m1_28490_22513# m1_28490_22513# m1_27462_21586#
+ vss nfet$3
Xpfet$5_10 vdd vdd m1_23486_21590# m1_23356_21786# pfet$5
Xpfet$6_9 vdd vdd m1_29087_15778# m1_26217_17714# pfet$6
Xpfet$10_2 vdd vdd m1_n789_25858# m1_326_24346# pfet$10
Xpfet$4_6 vdd vdd vdd m1_6339_19850# m1_8137_20152# m1_8137_20152# pfet$4
Xpfet$2_22 vdd vdd m1_3015_15778# m1_3372_16080# pfet$2
Xpfet$2_11 vdd vdd m1_9485_17714# m1_9944_16080# pfet$2
Xpfet$2_33 vdd vdd m1_5892_17518# m1_5302_17714# pfet$2
Xpfet$2_99 vdd m1_23109_16202# m1_22624_17518# m1_23007_17836# pfet$2
Xpfet$2_88 vdd vdd m1_18441_17518# m1_17851_17714# pfet$2
Xpfet$2_77 vdd vdd m1_17851_17714# m1_18310_16080# pfet$2
Xpfet$2_66 vdd vdd m1_24904_15778# m1_22034_17714# pfet$2
Xnfet$9_9 m1_n10452_25858# vss m1_27031_17343# vss nfet$9
Xpfet$2_3 vdd m1_11381_15778# m1_10560_16202# m1_10299_17343# pfet$2
Xpfet$2_44 vdd vdd m1_649_17714# m1_1119_17714# pfet$2
Xpfet$2_55 vdd vdd m1_n2474_17518# m1_n3064_17714# pfet$2
Xnfet$29_4 m1_n10572_23922# vss m1_n9952_24224# vss nfet$29
Xnfet$34_2 m1_n6839_21786# vss m1_n6973_21481# vss nfet$34
Xnfet$27_1 m1_n8283_19850# vss m1_n6856_24542# vss nfet$27
Xnfet$10_13 m1_32675_25947# vss m1_32817_25662# vss nfet$10
Xnfet$7_6 m1_9015_17714# vss m1_12935_19550# vss nfet$7
Xpfet$2_110 vdd vdd m1_10458_17836# m1_10299_17343# pfet$2
Xnfet$13_7 m1_34278_25658# m1_34278_25658# vss vss m1_34737_25502# vss nfet$13
Xnfet$6_16 m1_26873_21786# vss m1_27003_21590# vss nfet$6
Xnfet$21_23 m1_18926_16202# m1_18926_16202# vss vss m1_18408_16398# vss nfet$21
Xnfet$21_12 m1_n1168_15778# m1_n1168_15778# m1_n1278_18030# m1_n1278_18030# m1_n1042_17358#
+ vss nfet$21
Xpfet$26_0 vdd vdd m1_n4485_20152# m1_n3822_20130# pfet$26
Xnfet$5_3 m1_n7513_20152# vss m1_9944_16080# vss nfet$5
Xnfet$11_4 m1_32193_25858# m1_34278_25658# m1_35071_24542# vss nfet$11
Xpfet$12_6 vdd vdd m1_31535_19792# m1_14422_22513# pfet$12
Xnfet$3_17 m1_12935_21590# m1_12935_21590# m1_14422_22513# m1_14422_22513# m1_13394_21586#
+ vss nfet$3
Xnfet$3_0 m1_n1133_21590# m1_n1133_21590# m1_354_22513# m1_354_22513# m1_n674_21586#
+ vss nfet$3
Xpfet$5_11 vdd vdd m1_18705_21786# m1_18073_21786# pfet$5
Xpfet$10_3 vdd m1_n646_24542# vdd m1_326_24346# pfet$10
Xpfet$4_7 vdd vdd vdd m1_6975_19550# m1_965_15478# m1_965_15478# pfet$4
Xpfet$2_89 vdd vdd m1_22848_17343# m1_25747_17714# pfet$2
Xpfet$2_78 vdd vdd m1_13514_15478# sd4 pfet$2
Xpfet$2_67 vdd m1_22034_17714# vdd m1_23109_16202# pfet$2
Xpfet$2_12 vdd m1_3989_15778# m1_3372_16080# m1_2092_17836# pfet$2
Xpfet$2_4 vdd m1_9485_17714# vdd m1_10560_16202# pfet$2
Xpfet$2_23 vdd m1_5302_17714# vdd m1_6377_16202# pfet$2
Xpfet$2_34 vdd vdd m1_5761_16080# m1_n7513_20152# pfet$2
Xpfet$2_45 vdd vdd m1_9944_16080# m1_n7513_20152# pfet$2
Xpfet$2_56 vdd m1_n1278_18030# vdd m1_n2605_16080# pfet$2
Xnfet$29_5 m1_n10933_25858# vss m1_n10796_25662# vss nfet$29
Xnfet$7_7 m1_5148_15478# vss m1_11654_20152# vss nfet$7
Xnfet$6_17 m1_25107_21786# vss m1_25739_21786# vss nfet$6
Xpfet$2_100 vdd vdd m1_23820_18030# m1_23930_15778# pfet$2
Xnfet$21_24 m1_18310_16080# m1_18310_16080# m1_17851_17714# m1_17851_17714# m1_18408_16398#
+ vss nfet$21
Xnfet$21_13 m1_n2605_16080# m1_n2605_16080# vss vss m1_n1042_17358# vss nfet$21
Xpfet$19_0 vdd vdd m1_n7247_17714# m1_n6788_16080# pfet$19
Xpfet$26_1 vdd m1_n4485_21904# vdd m1_9624_19404# pfet$26
Xnfet$32_0 m1_n7186_25858# vss m1_n7320_25516# vss nfet$32
Xnfet$5_4 m1_10299_17343# m1_10560_16202# m1_10075_17518# vss nfet$5
Xpfet$12_7 vdd vdd m1_31535_22102# m1_354_22513# pfet$12
Xnfet$11_5 m1_32330_25662# m1_33174_24224# m1_34278_25658# vss nfet$11
Xnfet$3_1 m1_n1263_21786# m1_n1263_21786# m1_354_22513# m1_354_22513# m1_n42_21586#
+ vss nfet$3
Xpfet$5_12 vdd vdd m1_16452_21590# m1_16322_21786# pfet$5
Xpfet$10_4 vdd vdd m1_32675_25947# m1_33790_24346# pfet$10
Xpfet$4_8 vdd m1_9624_19404# m1_9624_19404# m1_10492_19550# m1_4832_17714# m1_4832_17714#
+ pfet$4
Xpfet$2_79 vdd m1_15564_15778# m1_14743_16202# m1_14482_17343# pfet$2
Xpfet$2_68 vdd vdd m1_22034_17714# m1_22493_16080# pfet$2
Xpfet$2_13 vdd vdd m1_5148_15478# sd6 pfet$2
Xpfet$2_24 vdd m1_6377_16202# m1_5892_17518# m1_6275_17836# pfet$2
Xpfet$2_35 vdd vdd m1_9015_17714# m1_9485_17714# pfet$2
Xpfet$2_46 vdd vdd m1_n2250_17343# m1_649_17714# pfet$2
Xpfet$2_57 vdd m1_n1989_16202# m1_n2474_17518# m1_n2091_17836# pfet$2
Xnfet$29_6 m1_n10452_25858# vss m1_n10309_25662# vss nfet$29
Xpfet$2_5 vdd m1_7198_15778# m1_6377_16202# m1_6116_17343# pfet$2
Xnfet$7_8 m1_n7383_17599# vss m1_n1133_19550# vss nfet$7
Xpfet$2_101 vdd vdd m1_19637_18030# m1_19747_15778# pfet$2
Xnfet$25_0 m1_n5351_15778# m1_n5351_15778# m1_n5461_18030# m1_n5461_18030# m1_n5225_17358#
+ vss nfet$25
Xpfet$19_1 vdd m1_n7247_17714# vdd m1_n6172_16202# pfet$19
Xpfet$26_2 vdd m1_n5227_21418# vdd m1_2590_19404# pfet$26
Xnfet$32_1 m1_n6856_24542# vss m1_n6111_25858# vss nfet$32
Xnfet$21_25 m1_14743_16202# m1_14743_16202# vss vss m1_14225_16398# vss nfet$21
Xnfet$5_5 m1_10458_17836# m1_11738_16080# m1_11271_18030# vss nfet$5
Xnfet$21_14 m1_n2605_16080# m1_n2605_16080# m1_n3064_17714# m1_n3064_17714# m1_n2507_16398#
+ vss nfet$21
Xnfet$11_6 m1_32193_25858# m1_32817_25662# m1_32554_23922# vss nfet$11
Xpfet$31_0 vdd vdd m1_n5227_20152# m1_n2543_20130# pfet$31
Xpfet$5_13 vdd vdd m1_15188_21786# m1_14556_21786# pfet$5
Xnfet$3_2 m1_9288_21786# m1_9288_21786# m1_9645_21447# m1_9645_21447# m1_10509_21586#
+ vss nfet$3
Xpfet$10_5 vdd m1_32675_25947# vdd m1_34278_25658# pfet$10
Xpfet$4_9 vdd m1_9624_19404# m1_9624_19404# m1_9856_19850# m1_9418_19550# m1_9418_19550#
+ pfet$4
Xpfet$2_69 vdd vdd m1_20721_15778# m1_17851_17714# pfet$2
Xpfet$2_14 vdd vdd m1_2092_17836# m1_1933_17343# pfet$2
Xpfet$2_25 vdd vdd m1_1709_17518# m1_1119_17714# pfet$2
Xpfet$2_36 vdd vdd m1_6116_17343# m1_9015_17714# pfet$2
Xpfet$2_47 vdd m1_11738_16080# m1_11271_18030# m1_10299_17343# pfet$2
Xpfet$2_58 vdd vdd m1_n3534_17714# m1_n3064_17714# pfet$2
Xnfet$29_7 m1_n7320_25516# vss m1_n2567_23922# vss nfet$29
Xpfet$2_6 vdd vdd m1_7198_15778# m1_7555_16080# pfet$2
Xnfet$7_9 m1_25747_17714# vss m1_27003_19550# vss nfet$7
Xpfet$2_102 vdd vdd m1_13198_17714# m1_13668_17714# pfet$2
Xpfet$19_2 vdd vdd m1_n5461_18030# m1_n5351_15778# pfet$19
Xpfet$26_3 vdd vdd m1_n5227_21418# m1_6107_19404# pfet$26
Xnfet$21_26 m1_14127_16080# m1_14127_16080# m1_13668_17714# m1_13668_17714# m1_14225_16398#
+ vss nfet$21
Xnfet$18_0 m1_34093_19792# vss m1_34843_21786# vss nfet$18
Xnfet$5_6 m1_6116_17343# vss m1_6275_17836# vss nfet$5
Xnfet$25_1 m1_n6788_16080# m1_n6788_16080# vss vss m1_n5225_17358# vss nfet$25
Xnfet$21_15 m1_n1989_16202# m1_n1989_16202# vss vss m1_n2507_16398# vss nfet$21
Xnfet$11_7 m1_32330_25662# m1_32554_23922# m1_32818_24542# vss nfet$11
Xpfet$31_1 vdd m1_n4485_20152# vdd m1_n3206_20274# pfet$31
Xpfet$24_0 vdd vdd m1_n7320_25516# m1_n7186_25858# pfet$24
Xnfet$3_3 m1_9418_21590# m1_9418_21590# m1_9645_21447# m1_9645_21447# m1_9877_21586#
+ vss nfet$3
Xpfet$10_6 vdd vdd m1_32818_24542# m1_33174_24224# pfet$10
Xpfet$5_14 vdd vdd m1_19969_21590# m1_19839_21786# pfet$5
Xnfet$1_0 m1_4509_24346# m1_4509_24346# vss vss m1_3991_24542# vss nfet$1
Xpfet$9_0 vdd vdd m1_n647_25662# m1_n789_25858# pfet$9
Xpfet$2_15 vdd vdd m1_5302_17714# m1_5761_16080# pfet$2
Xpfet$2_26 vdd vdd m1_4832_17714# m1_5302_17714# pfet$2
Xpfet$2_37 vdd m1_7555_16080# m1_7088_18030# m1_6116_17343# pfet$2
Xpfet$2_48 vdd vdd m1_n3064_17714# m1_n2605_16080# pfet$2
Xpfet$2_59 vdd vdd m1_n2605_16080# m1_n7513_20152# pfet$2
Xnfet$29_8 m1_n4623_25487# vss m1_n4464_25980# vss nfet$29
Xpfet$2_7 vdd vdd m1_6275_17836# m1_6116_17343# pfet$2
Xnfet$1_20 m1_21241_24346# m1_21241_24346# m1_20126_25858# m1_20126_25858# m1_22188_25502#
+ vss nfet$1
Xpfet$2_103 vdd m1_14743_16202# m1_14258_17518# m1_14641_17836# pfet$2
Xnfet$21_27 m1_18310_16080# m1_18310_16080# vss vss m1_19873_17358# vss nfet$21
Xnfet$21_16 m1_19747_15778# m1_19747_15778# m1_19637_18030# m1_19637_18030# m1_19873_17358#
+ vss nfet$21
Xnfet$18_1 m1_30256_19792# vss m1_32818_20470# vss nfet$18
Xnfet$5_7 m1_9485_17714# vss m1_10075_17518# vss nfet$5
Xnfet$25_2 m1_n6788_16080# m1_n6788_16080# m1_n7247_17714# m1_n7247_17714# m1_n6690_16398#
+ vss nfet$25
Xpfet$19_3 vdd m1_n5461_18030# vdd m1_n6788_16080# pfet$19
Xpfet$26_4 vdd vdd m1_n4485_21904# m1_n3822_21786# pfet$26
Xpfet$17_0 vdd vdd fout m1_34093_22102# pfet$17
Xpfet$31_2 vdd m1_n5227_20152# vdd m1_n1927_20274# pfet$31
Xnfet$30_0 m1_n9952_24224# m1_n9952_24224# m1_n10308_24542# m1_n10308_24542# m1_n9854_24542#
+ vss nfet$30
Xpfet$24_1 vdd vdd m1_n6111_25858# m1_n6856_24542# pfet$24
Xnfet$3_4 m1_5901_21590# m1_5901_21590# m1_7388_22513# m1_7388_22513# m1_6360_21586#
+ vss nfet$3
Xpfet$10_7 vdd m1_32818_24542# vdd m1_33790_24346# pfet$10
Xpfet$5_15 vdd vdd m1_27003_21590# m1_26873_21786# pfet$5
Xnfet$1_1 m1_3893_24224# m1_3893_24224# m1_3537_24542# m1_3537_24542# m1_3991_24542#
+ vss nfet$1
Xpfet$9_1 vdd vdd m1_n1134_25662# m1_n1271_25858# pfet$9
Xpfet$2_16 vdd vdd m1_3989_15778# m1_1119_17714# pfet$2
Xpfet$2_27 vdd m1_2194_16202# m1_1709_17518# m1_2092_17836# pfet$2
Xpfet$2_38 vdd vdd m1_7088_18030# m1_7198_15778# pfet$2
Xpfet$2_49 vdd m1_n194_15778# m1_n811_16080# m1_n2091_17836# pfet$2
Xpfet$2_8 vdd vdd m1_9331_15478# sd5 pfet$2
Xnfet$29_9 m1_n3184_24224# vss m1_n3541_23922# vss nfet$29
Xnfet$1_21 m1_28991_24224# m1_28991_24224# m1_28635_24542# m1_28635_24542# m1_29089_24542#
+ vss nfet$1
Xnfet$1_10 m1_17546_25658# m1_17546_25658# vss vss m1_18005_25502# vss nfet$1
Xpfet$2_104 vdd vdd m1_14127_16080# m1_n7513_20152# pfet$2
Xnfet$21_17 m1_22493_16080# m1_22493_16080# vss vss m1_24056_17358# vss nfet$21
Xnfet$18_2 m1_31535_19792# m1_32818_20470# vss vss nfet$18
Xpfet$19_4 vdd vdd m1_26217_17714# m1_26676_16080# pfet$19
Xnfet$25_3 m1_n6172_16202# m1_n6172_16202# vss vss m1_n6690_16398# vss nfet$25
Xpfet$26_5 vdd m1_n6839_21786# vdd m1_n5764_21786# pfet$26
Xnfet$5_8 m1_7555_16080# vss m1_7198_15778# vss nfet$5
Xpfet$31_3 vdd m1_n6839_20152# vdd m1_n927_19404# pfet$31
Xnfet$23_0 m1_35837_22102# vss m1_n7513_20152# vss nfet$23
Xnfet$30_1 m1_n9336_24346# m1_n9336_24346# m1_n8625_26174# m1_n8625_26174# m1_n8389_25502#
+ vss nfet$30
Xnfet$3_5 m1_2254_21786# m1_2254_21786# m1_3871_22513# m1_3871_22513# m1_3475_21586#
+ vss nfet$3
Xpfet$5_16 vdd vdd m1_29256_21786# m1_28624_21786# pfet$5
Xnfet$1_2 m1_4997_25658# m1_4997_25658# vss vss m1_5456_25502# vss nfet$1
Xnfet$4_10 m1_9015_17714# m1_9015_17714# vss vss m1_14005_20470# vss nfet$4
Xpfet$9_2 vdd vdd m1_n1271_25858# m1_n10452_25858# pfet$9
Xpfet$2_17 vdd vdd m1_n2091_17836# m1_n2250_17343# pfet$2
Xpfet$2_9 vdd vdd m1_8172_15778# m1_5302_17714# pfet$2
Xpfet$2_28 vdd m1_2905_18030# vdd m1_1578_16080# pfet$2
Xpfet$2_39 vdd m1_7088_18030# vdd m1_5761_16080# pfet$2
Xnfet$1_22 m1_29607_24346# m1_29607_24346# vss vss m1_29089_24542# vss nfet$1
Xnfet$1_11 m1_16442_24224# m1_16442_24224# m1_16086_24542# m1_16086_24542# m1_16540_24542#
+ vss nfet$1
Xpfet$2_105 vdd vdd m1_14258_17518# m1_13668_17714# pfet$2
Xnfet$18_3 m1_30256_22102# vss m1_32818_21586# vss nfet$18
Xnfet$21_18 m1_23930_15778# m1_23930_15778# m1_23820_18030# m1_23820_18030# m1_24056_17358#
+ vss nfet$21
Xnfet$25_4 m1_28113_15778# m1_28113_15778# m1_28003_18030# m1_28003_18030# m1_28239_17358#
+ vss nfet$25
Xpfet$19_5 vdd m1_26217_17714# vdd m1_27292_16202# pfet$19
Xpfet$26_6 vdd vdd m1_n6973_21481# m1_n6839_21786# pfet$26
Xnfet$5_9 sd5 vss m1_9331_15478# vss nfet$5
Xnfet$7_10 m1_26063_15478# vss m1_29239_20152# vss nfet$7
Xnfet$16_0 m1_34843_21786# m1_34843_21786# m1_34093_22102# m1_34093_22102# m1_34329_21430#
+ vss nfet$16
Xpfet$31_4 vdd vdd m1_n6839_20152# m1_n6973_21481# pfet$31
Xnfet$30_2 m1_n8848_25658# m1_n8848_25658# vss vss m1_n8389_25502# vss nfet$30
Xnfet$3_6 m1_2384_21590# m1_2384_21590# m1_3871_22513# m1_3871_22513# m1_2843_21586#
+ vss nfet$3
Xpfet$5_17 vdd vdd m1_25739_21786# m1_25107_21786# pfet$5
Xpfet$22_0 vdd vdd vdd m1_n6624_23622# m1_n7082_23622# m1_n7082_23622# pfet$22
Xnfet$1_3 m1_4509_24346# m1_4509_24346# m1_3394_25858# m1_3394_25858# m1_5456_25502#
+ vss nfet$1
Xnfet$4_11 m1_13198_17714# m1_13198_17714# vss vss m1_17522_20470# vss nfet$4
Xpfet$9_3 vdd vdd m1_1607_24542# m1_n789_25858# pfet$9
Xpfet$2_18 vdd m1_1119_17714# vdd m1_2194_16202# pfet$2
Xpfet$2_29 vdd vdd m1_1578_16080# m1_n7513_20152# pfet$2
Xpfet$7_0 vdd vdd m1_2384_19550# m1_n3534_17714# pfet$7
Xnfet$1_23 m1_25424_24346# m1_25424_24346# m1_24309_25858# m1_24309_25858# m1_26371_25502#
+ vss nfet$1
Xnfet$1_12 m1_17058_24346# m1_17058_24346# m1_15943_25858# m1_15943_25858# m1_18005_25502#
+ vss nfet$1
Xpfet$2_106 vdd vdd m1_14482_17343# m1_17381_17714# pfet$2
Xpfet$19_6 vdd vdd m1_28003_18030# m1_28113_15778# pfet$19
Xnfet$25_5 m1_26676_16080# m1_26676_16080# vss vss m1_28239_17358# vss nfet$25
Xpfet$26_7 vdd vdd m1_n6839_21786# m1_n6380_21786# pfet$26
Xnfet$21_19 m1_23109_16202# m1_23109_16202# vss vss m1_22591_16398# vss nfet$21
Xnfet$16_1 m1_28490_22513# m1_28490_22513# vss vss m1_34329_21430# vss nfet$16
Xnfet$7_11 m1_9331_15478# vss m1_15171_20152# vss nfet$7
Xnfet$30_3 m1_n9336_24346# m1_n9336_24346# vss vss m1_n9854_24542# vss nfet$30
Xnfet$3_7 m1_5771_21786# m1_5771_21786# m1_7388_22513# m1_7388_22513# m1_6992_21586#
+ vss nfet$3
Xpfet$15_0 vdd m1_34093_22102# vdd m1_28490_22513# pfet$15
Xnfet$1_4 m1_12259_24224# m1_12259_24224# m1_11903_24542# m1_11903_24542# m1_12357_24542#
+ vss nfet$1
Xpfet$22_1 vdd m1_n6856_24542# m1_n6856_24542# m1_n6624_23622# m1_n8283_19850# m1_n8283_19850#
+ pfet$22
Xnfet$4_12 m1_16452_19550# m1_16452_19550# vss vss m1_16890_20470# vss nfet$4
Xpfet$9_4 vdd vdd m1_488_21786# m1_n789_25858# pfet$9
Xpfet$2_19 vdd m1_3015_15778# m1_2194_16202# m1_1933_17343# pfet$2
Xpfet$7_1 vdd vdd m1_4620_20152# m1_n3218_15478# pfet$7
Xnfet$1_24 m1_30095_25658# m1_30095_25658# vss vss m1_30554_25502# vss nfet$1
Xnfet$1_13 m1_13363_25658# m1_13363_25658# vss vss m1_13822_25502# vss nfet$1
Xpfet$2_107 vdd m1_15921_16080# m1_15454_18030# m1_14482_17343# pfet$2
Xpfet$19_7 vdd m1_28003_18030# vdd m1_26676_16080# pfet$19
Xnfet$25_6 m1_27292_16202# m1_27292_16202# vss vss m1_26774_16398# vss nfet$25
Xnfet$16_2 m1_9645_21447# m1_9645_21447# vss vss m1_30492_21430# vss nfet$16
Xnfet$7_12 m1_13514_15478# vss m1_18688_20152# vss nfet$7
Xnfet$30_4 m1_n4978_24224# m1_n4978_24224# m1_n10452_25858# m1_n10452_25858# m1_n4880_24542#
+ vss nfet$30
Xnfet$3_8 m1_23486_21590# m1_23486_21590# m1_24973_22513# m1_24973_22513# m1_23945_21586#
+ vss nfet$3
Xpfet$15_1 vdd vdd m1_34093_22102# m1_34843_21786# pfet$15
Xnfet$1_5 m1_8692_24346# m1_8692_24346# vss vss m1_8174_24542# vss nfet$1
Xnfet$21_0 m1_7198_15778# m1_7198_15778# m1_7088_18030# m1_7088_18030# m1_7324_17358#
+ vss nfet$21
Xnfet$4_13 m1_19969_19550# m1_19969_19550# vss vss m1_20407_20470# vss nfet$4
Xpfet$9_5 vdd vdd m1_326_24346# m1_n7513_20152# pfet$9
Xpfet$7_2 vdd vdd m1_1103_20152# m1_n7401_15478# pfet$7
Xnfet$1_25 m1_29607_24346# m1_29607_24346# m1_28492_25858# m1_28492_25858# m1_30554_25502#
+ vss nfet$1
Xnfet$1_14 m1_12875_24346# m1_12875_24346# m1_11760_25858# m1_11760_25858# m1_13822_25502#
+ vss nfet$1
Xpfet$3_30 vdd vdd vdd m1_17539_22402# m1_16322_21786# m1_16322_21786# pfet$3
Xpfet$2_108 vdd vdd m1_15454_18030# m1_15564_15778# pfet$2
Xnfet$25_7 m1_26676_16080# m1_26676_16080# m1_26217_17714# m1_26217_17714# m1_26774_16398#
+ vss nfet$25
Xnfet$7_13 m1_13198_17714# vss m1_16452_19550# vss nfet$7
Xnfet$30_5 m1_n4362_24346# m1_n4362_24346# vss vss m1_n4880_24542# vss nfet$30
Xnfet$16_3 m1_7388_22513# m1_7388_22513# m1_30256_22102# m1_30256_22102# m1_30492_21430#
+ vss nfet$16
Xnfet$3_9 m1_23356_21786# m1_23356_21786# m1_24973_22513# m1_24973_22513# m1_24577_21586#
+ vss nfet$3
Xpfet$15_2 vdd vdd m1_30256_22102# m1_7388_22513# pfet$15
Xnfet$21_1 m1_5761_16080# m1_5761_16080# vss vss m1_7324_17358# vss nfet$21
Xnfet$14_0 m1_11039_21786# m1_11039_21786# vss vss m1_9877_21586# vss nfet$14
Xnfet$1_6 m1_8076_24224# m1_8076_24224# m1_7720_24542# m1_7720_24542# m1_8174_24542#
+ vss nfet$1
Xnfet$4_14 m1_17381_17714# m1_17381_17714# vss vss m1_21039_20470# vss nfet$4
Xpfet$9_6 vdd vdd m1_n290_24224# m1_n910_23922# pfet$9
Xpfet$20_0 vdd m1_n4377_15778# m1_n4994_16080# m1_n6274_17836# pfet$20
Xnfet$14_10 m1_21590_21786# m1_21590_21786# vss vss m1_20428_21586# vss nfet$14
Xpfet$7_3 vdd vdd m1_5901_19550# m1_649_17714# pfet$7
Xnfet$1_26 m1_25912_25658# m1_25912_25658# vss vss m1_26371_25502# vss nfet$1
Xnfet$1_15 m1_25424_24346# m1_25424_24346# vss vss m1_24906_24542# vss nfet$1
Xpfet$3_31 vdd vdd vdd m1_27462_22102# m1_27003_21590# m1_27003_21590# pfet$3
Xpfet$3_20 vdd vdd vdd m1_20428_22102# m1_19969_21590# m1_19969_21590# pfet$3
Xpfet$2_109 vdd vdd m1_10299_17343# m1_13198_17714# pfet$2
Xpfet$5_0 vdd vdd m1_n1133_21590# m1_n1263_21786# pfet$5
Xnfet$2_80 m1_28147_25662# m1_28991_24224# m1_30095_25658# vss nfet$2
Xnfet$7_14 m1_21564_17714# vss m1_23486_19550# vss nfet$7
Xnfet$30_6 m1_n4978_24224# m1_n4978_24224# vss vss m1_n3415_25502# vss nfet$30
Xnfet$22_10 m1_9331_15478# m1_9331_15478# m1_n3822_21786# m1_n3822_21786# m1_13373_20470#
+ vss nfet$22
Xnfet$8_0 sd9 vss m1_n7401_15478# vss nfet$8
Xpfet$15_3 vdd m1_31535_22102# vdd m1_3871_22513# pfet$15
Xnfet$21_2 m1_9944_16080# m1_9944_16080# vss vss m1_11507_17358# vss nfet$21
Xnfet$14_1 m1_11671_21786# m1_11671_21786# vss vss m1_10509_21586# vss nfet$14
Xnfet$1_7 m1_9180_25658# m1_9180_25658# vss vss m1_9639_25502# vss nfet$1
Xnfet$4_15 m1_21564_17714# m1_21564_17714# vss vss m1_24556_20470# vss nfet$4
Xpfet$9_7 vdd vdd m1_32330_25662# m1_32193_25858# pfet$9
Xpfet$20_1 vdd m1_n5351_15778# m1_n6172_16202# m1_n6433_17343# pfet$20
Xpfet$13_0 vdd m1_n647_25662# m1_n910_23922# m1_n1134_25662# pfet$13
Xpfet$7_4 vdd vdd m1_12935_19550# m1_9015_17714# pfet$7
Xnfet$14_11 m1_22222_21786# m1_22222_21786# vss vss m1_21060_21586# vss nfet$14
Xnfet$5_80 m1_18824_17836# m1_19747_15778# m1_18926_16202# vss nfet$5
Xnfet$1_27 m1_12875_24346# m1_12875_24346# vss vss m1_12357_24542# vss nfet$1
Xpfet$3_32 vdd m1_28490_22513# m1_28490_22513# m1_28090_22402# m1_28624_21786# m1_28624_21786#
+ pfet$3
Xnfet$1_16 m1_24808_24224# m1_24808_24224# m1_24452_24542# m1_24452_24542# m1_24906_24542#
+ vss nfet$1
Xpfet$3_21 vdd vdd vdd m1_21056_22402# m1_19839_21786# m1_19839_21786# pfet$3
Xpfet$3_10 vdd m1_3871_22513# m1_3871_22513# m1_2843_22102# m1_4637_21786# m1_4637_21786#
+ pfet$3
Xpfet$5_1 vdd vdd m1_11671_21786# m1_11039_21786# pfet$5
Xpfet$1_110 vdd m1_11903_24542# vdd m1_12875_24346# pfet$1
Xnfet$2_81 m1_n7513_20152# vss m1_25424_24346# vss nfet$2
Xnfet$2_70 m1_21590_21786# vss m1_28010_25858# vss nfet$2
Xnfet$37_0 m1_n6839_20152# vss m1_n8145_21908# vss nfet$37
Xnfet$7_15 m1_17697_15478# vss m1_22205_20152# vss nfet$7
Xnfet$30_7 m1_n3541_23922# m1_n3541_23922# m1_n3651_26174# m1_n3651_26174# m1_n3415_25502#
+ vss nfet$30
Xnfet$22_11 m1_15171_20152# m1_15171_20152# m1_n3822_21786# m1_n3822_21786# m1_14005_20470#
+ vss nfet$22
Xnfet$8_1 sd2 vss m1_21880_15478# vss nfet$8
Xpfet$15_4 vdd m1_30256_22102# vdd m1_9645_21447# pfet$15
Xnfet$1_8 m1_8692_24346# m1_8692_24346# m1_7577_25858# m1_7577_25858# m1_9639_25502#
+ vss nfet$1
Xnfet$21_3 m1_11381_15778# m1_11381_15778# m1_11271_18030# m1_11271_18030# m1_11507_17358#
+ vss nfet$21
Xnfet$14_2 m1_8154_21786# m1_8154_21786# vss vss m1_6992_21586# vss nfet$14
Xnfet$4_16 m1_23486_19550# m1_23486_19550# vss vss m1_23924_20470# vss nfet$4
Xpfet$9_8 vdd vdd m1_33174_24224# m1_32554_23922# pfet$9
Xpfet$6_10 vdd vdd m1_27031_17343# m1_n10452_25858# pfet$6
Xpfet$20_2 vdd m1_n4994_16080# m1_n5461_18030# m1_n6433_17343# pfet$20
Xpfet$13_1 vdd m1_n910_23922# m1_n646_24542# m1_n1271_25858# pfet$13
Xpfet$7_5 vdd vdd m1_8137_20152# m1_965_15478# pfet$7
Xnfet$5_81 m1_13198_17714# vss m1_10299_17343# vss nfet$5
Xnfet$14_12 m1_18073_21786# m1_18073_21786# vss vss m1_16911_21586# vss nfet$14
Xnfet$5_70 m1_n7513_20152# vss m1_18310_16080# vss nfet$5
Xpfet$3_33 vdd m1_28490_22513# m1_28490_22513# m1_27462_22102# m1_29256_21786# m1_29256_21786#
+ pfet$3
Xnfet$1_17 m1_20625_24224# m1_20625_24224# m1_20269_24542# m1_20269_24542# m1_20723_24542#
+ vss nfet$1
Xpfet$3_22 vdd m1_21456_22513# m1_21456_22513# m1_20428_22102# m1_22222_21786# m1_22222_21786#
+ pfet$3
Xpfet$3_11 vdd vdd vdd m1_2843_22102# m1_2384_21590# m1_2384_21590# pfet$3
Xpfet$5_2 vdd vdd m1_12935_21590# m1_12805_21786# pfet$5
Xpfet$1_100 vdd vdd m1_29607_24346# m1_n7513_20152# pfet$1
Xnfet$2_82 m1_11415_25662# m1_12259_24224# m1_13363_25658# vss nfet$2
Xnfet$2_71 m1_28147_25662# m1_28371_23922# m1_28635_24542# vss nfet$2
Xnfet$2_60 pd6 vss m1_16322_21786# vss nfet$2
Xpfet$9_10 vdd vdd m1_35071_24542# m1_32675_25947# pfet$9
Xnfet$7_16 m1_17381_17714# vss m1_19969_19550# vss nfet$7
Xnfet$8_2 sd1 vss m1_26063_15478# vss nfet$8
Xnfet$22_12 m1_18688_20152# m1_18688_20152# m1_n1927_20274# m1_n1927_20274# m1_17522_20470#
+ vss nfet$22
Xnfet$1_9 m1_17058_24346# m1_17058_24346# vss vss m1_16540_24542# vss nfet$1
Xnfet$21_4 m1_10560_16202# m1_10560_16202# vss vss m1_10042_16398# vss nfet$21
Xnfet$14_3 m1_7522_21786# m1_7522_21786# vss vss m1_6360_21586# vss nfet$14
Xnfet$4_17 m1_12935_19550# m1_12935_19550# vss vss m1_13373_20470# vss nfet$4
Xpfet$9_9 vdd vdd m1_28624_21786# m1_32675_25947# pfet$9
Xpfet$6_11 vdd vdd m1_26807_17518# m1_26217_17714# pfet$6
Xnfet$12_0 pd1 vss m1_n1263_21786# vss nfet$12
Xpfet$20_3 vdd m1_n6172_16202# m1_n6657_17518# m1_n6274_17836# pfet$20
Xpfet$13_2 vdd m1_n290_24224# m1_814_25658# m1_n1271_25858# pfet$13
Xnfet$5_82 m1_10299_17343# vss m1_10458_17836# vss nfet$5
Xnfet$14_13 m1_18705_21786# m1_18705_21786# vss vss m1_17543_21586# vss nfet$14
Xnfet$5_71 m1_14641_17836# m1_15921_16080# m1_15454_18030# vss nfet$5
Xnfet$5_60 m1_18665_17343# vss m1_18824_17836# vss nfet$5
Xpfet$7_6 vdd vdd m1_9418_19550# m1_4832_17714# pfet$7
Xnfet$1_18 m1_21241_24346# m1_21241_24346# vss vss m1_20723_24542# vss nfet$1
Xpfet$3_12 vdd vdd vdd m1_3471_22402# m1_2254_21786# m1_2254_21786# pfet$3
Xpfet$3_34 vdd vdd vdd m1_28090_22402# m1_26873_21786# m1_26873_21786# pfet$3
Xpfet$3_23 vdd vdd vdd m1_23945_22102# m1_23486_21590# m1_23486_21590# pfet$3
Xpfet$5_3 vdd vdd m1_9418_21590# m1_9288_21786# pfet$5
Xpfet$1_101 vdd vdd m1_28010_25858# m1_21590_21786# pfet$1
Xnfet$2_72 m1_23827_25858# m1_25912_25658# m1_26705_24542# vss nfet$2
Xnfet$2_61 m1_23964_25662# m1_24808_24224# m1_25912_25658# vss nfet$2
Xnfet$2_50 m1_n7513_20152# vss m1_21241_24346# vss nfet$2
Xpfet$3_0 vdd vdd vdd m1_n674_22102# m1_n1133_21590# m1_n1133_21590# pfet$3
Xnfet$7_17 m1_21880_15478# vss m1_25722_20152# vss nfet$7
Xpfet$9_11 vdd vdd m1_32817_25662# m1_32675_25947# pfet$9
Xnfet$22_13 m1_13514_15478# m1_13514_15478# m1_n1927_20274# m1_n1927_20274# m1_16890_20470#
+ vss nfet$22
Xpfet$29_0 vdd vdd vdd m1_n8047_19550# m1_n7513_20152# m1_n7513_20152# pfet$29
Xnfet$21_5 m1_9944_16080# m1_9944_16080# m1_9485_17714# m1_9485_17714# m1_10042_16398#
+ vss nfet$21
Xnfet$14_4 m1_1120_21786# m1_1120_21786# vss vss m1_n42_21586# vss nfet$14
Xnfet$6_0 m1_n1263_21786# vss m1_n1133_21590# vss nfet$6
Xpfet$6_12 vdd vdd m1_26676_16080# m1_n7513_20152# pfet$6
Xpfet$20_4 vdd m1_28113_15778# m1_27292_16202# m1_27031_17343# pfet$20
Xpfet$13_3 vdd m1_814_25658# m1_1607_24542# m1_n1134_25662# pfet$13
Xnfet$12_1 pd2 vss m1_2254_21786# vss nfet$12
Xpfet$11_0 vdd vdd vdd m1_33050_22344# m1_31535_22102# m1_31535_22102# pfet$11
Xnfet$14_14 m1_15188_21786# m1_15188_21786# vss vss m1_14026_21586# vss nfet$14
Xnfet$5_72 m1_17851_17714# vss m1_18441_17518# vss nfet$5
Xnfet$5_61 m1_20104_16080# vss m1_19747_15778# vss nfet$5
Xnfet$5_50 m1_25747_17714# vss m1_22848_17343# vss nfet$5
Xpfet$7_7 vdd vdd m1_11654_20152# m1_5148_15478# pfet$7
Xnfet$1_19 m1_21729_25658# m1_21729_25658# vss vss m1_22188_25502# vss nfet$1
Xpfet$27_10 vdd vdd m1_n10933_25858# fin pfet$27
Xpfet$3_35 vdd vdd vdd m1_13394_22102# m1_12935_21590# m1_12935_21590# pfet$3
Xpfet$3_24 vdd m1_17939_22513# m1_17939_22513# m1_16911_22102# m1_18705_21786# m1_18705_21786#
+ pfet$3
Xpfet$3_13 vdd vdd vdd m1_6988_22402# m1_5771_21786# m1_5771_21786# pfet$3
Xpfet$5_4 vdd vdd m1_8154_21786# m1_7522_21786# pfet$5
Xpfet$1_102 vdd m1_28371_23922# m1_28635_24542# m1_28010_25858# pfet$1
Xnfet$2_73 m1_24309_25858# vss m1_21590_21786# vss nfet$2
Xnfet$2_62 m1_24188_23922# vss m1_24808_24224# vss nfet$2
Xnfet$2_51 m1_19644_25858# m1_21729_25658# m1_22522_24542# vss nfet$2
Xnfet$2_40 m1_15598_25662# m1_16442_24224# m1_17546_25658# vss nfet$2
Xpfet$3_1 vdd m1_7388_22513# m1_7388_22513# m1_6988_22402# m1_7522_21786# m1_7522_21786#
+ pfet$3
Xpfet$9_12 vdd vdd m1_32193_25858# m1_25107_21786# pfet$9
Xnfet$22_14 m1_22205_20152# m1_22205_20152# m1_n2543_20130# m1_n2543_20130# m1_21039_20470#
+ vss nfet$22
Xpfet$29_1 vdd m1_n8283_19850# m1_n8283_19850# m1_n8047_19550# m1_n8283_20611# m1_n8283_20611#
+ pfet$29
Xnfet$35_0 m1_n927_19404# m1_n927_19404# vss vss m1_n6282_20470# vss nfet$35
Xnfet$21_6 m1_1578_16080# m1_1578_16080# vss vss m1_3141_17358# vss nfet$21
Xnfet$14_5 m1_4005_21786# m1_4005_21786# vss vss m1_2843_21586# vss nfet$14
Xpfet$1_90 vdd vdd m1_24309_25858# m1_25424_24346# pfet$1
Xpfet$6_13 vdd vdd m1_25747_17714# m1_26217_17714# pfet$6
Xnfet$6_1 m1_11039_21786# vss m1_11671_21786# vss nfet$6
Xnfet$12_2 pd9 vss m1_26873_21786# vss nfet$12
Xpfet$13_4 vdd m1_33174_24224# m1_34278_25658# m1_32193_25858# pfet$13
Xpfet$20_5 vdd m1_29087_15778# m1_28470_16080# m1_27190_17836# pfet$20
Xnfet$14_15 m1_14556_21786# m1_14556_21786# vss vss m1_13394_21586# vss nfet$14
Xnfet$5_73 m1_13668_17714# vss m1_16538_15778# vss nfet$5
Xnfet$5_62 m1_18665_17343# m1_20721_15778# m1_20104_16080# vss nfet$5
Xnfet$5_51 m1_n7513_20152# vss m1_22493_16080# vss nfet$5
Xnfet$5_40 m1_n2250_17343# m1_n194_15778# m1_n811_16080# vss nfet$5
Xpfet$7_8 vdd vdd m1_n1133_19550# m1_n7383_17599# pfet$7
Xpfet$3_25 vdd m1_17939_22513# m1_17939_22513# m1_17539_22402# m1_18073_21786# m1_18073_21786#
+ pfet$3
Xpfet$3_14 vdd vdd vdd m1_n46_22402# m1_n1263_21786# m1_n1263_21786# pfet$3
Xpfet$27_11 vdd vdd m1_n9336_24346# vss pfet$27
Xpfet$5_5 vdd vdd m1_1120_21786# m1_488_21786# pfet$5
Xpfet$1_103 vdd vdd m1_28635_24542# m1_28991_24224# pfet$1
Xnfet$2_74 pd8 vss m1_23356_21786# vss nfet$2
Xnfet$2_63 m1_14556_21786# vss m1_19644_25858# vss nfet$2
Xnfet$2_52 m1_20126_25858# vss m1_22522_24542# vss nfet$2
Xnfet$2_41 pd5 vss m1_12805_21786# vss nfet$2
Xnfet$2_30 m1_n7513_20152# vss m1_17058_24346# vss nfet$2
Xpfet$3_2 vdd m1_7388_22513# m1_7388_22513# m1_6360_22102# m1_8154_21786# m1_8154_21786#
+ pfet$3
Xpfet$9_13 vdd vdd m1_33790_24346# m1_n7513_20152# pfet$9
Xnfet$35_1 m1_n2543_20130# m1_n2543_20130# m1_n5227_20152# m1_n5227_20152# m1_n2445_20470#
+ vss nfet$35
Xpfet$29_2 vdd m1_n8283_20611# m1_n8283_20611# m1_n8047_22344# m1_n8145_21908# m1_n8145_21908#
+ pfet$29
Xnfet$22_15 m1_17697_15478# m1_17697_15478# m1_n2543_20130# m1_n2543_20130# m1_20407_20470#
+ vss nfet$22
Xnfet$28_0 m1_n3822_20130# m1_n3822_20130# m1_n4485_20152# m1_n4485_20152# m1_n3724_20470#
+ vss nfet$28
Xnfet$21_7 m1_5761_16080# m1_5761_16080# m1_5302_17714# m1_5302_17714# m1_5859_16398#
+ vss nfet$21
Xnfet$14_6 m1_4637_21786# m1_4637_21786# vss vss m1_3475_21586# vss nfet$14
Xpfet$1_91 vdd vdd m1_23356_21786# pd8 pfet$1
Xpfet$1_80 vdd vdd m1_17058_24346# m1_n7513_20152# pfet$1
Xnfet$6_2 m1_12805_21786# vss m1_12935_21590# vss nfet$6
Xpfet$13_5 vdd m1_32817_25662# m1_32554_23922# m1_32330_25662# pfet$13
Xpfet$20_6 vdd m1_28470_16080# m1_28003_18030# m1_27031_17343# pfet$20
Xnfet$5_74 m1_14482_17343# vss m1_14641_17836# vss nfet$5
Xnfet$5_63 m1_13668_17714# vss m1_14258_17518# vss nfet$5
Xnfet$5_52 m1_23007_17836# m1_24287_16080# m1_23820_18030# vss nfet$5
Xpfet$7_9 vdd vdd m1_27003_19550# m1_25747_17714# pfet$7
Xnfet$5_30 sd6 vss m1_5148_15478# vss nfet$5
Xnfet$5_41 m1_n2091_17836# m1_n1168_15778# m1_n1989_16202# vss nfet$5
Xnfet$14_16 m1_28624_21786# m1_28624_21786# vss vss m1_27462_21586# vss nfet$14
Xnfet$10_0 m1_n10452_25858# vss m1_n1271_25858# vss nfet$10
Xpfet$3_26 vdd vdd vdd m1_16911_22102# m1_16452_21590# m1_16452_21590# pfet$3
Xpfet$3_15 vdd m1_354_22513# m1_354_22513# m1_n46_22402# m1_488_21786# m1_488_21786#
+ pfet$3
Xpfet$27_12 vdd vdd m1_n7082_23622# m1_n8625_26174# pfet$27
Xpfet$5_6 vdd vdd m1_5901_21590# m1_5771_21786# pfet$5
Xpfet$1_104 vdd m1_25912_25658# m1_26705_24542# m1_23964_25662# pfet$1
Xnfet$2_75 m1_28371_23922# vss m1_28991_24224# vss nfet$2
Xnfet$2_64 m1_19644_25858# vss m1_19781_25662# vss nfet$2
Xnfet$2_53 m1_23827_25858# m1_24451_25662# m1_24188_23922# vss nfet$2
Xnfet$2_42 m1_15943_25858# vss m1_16085_25662# vss nfet$2
Xnfet$2_31 m1_15943_25858# vss m1_18339_24542# vss nfet$2
Xnfet$2_20 pd3 vss m1_5771_21786# vss nfet$2
Xpfet$3_3 vdd m1_9645_21447# m1_9645_21447# m1_10505_22402# m1_11039_21786# m1_11039_21786#
+ pfet$3
Xnfet$22_16 m1_25722_20152# m1_25722_20152# m1_n3206_20274# m1_n3206_20274# m1_24556_20470#
+ vss nfet$22
Xnfet$28_1 m1_n1927_20274# m1_n1927_20274# vss vss m1_n2445_20470# vss nfet$28
Xpfet$29_3 vdd vdd vdd m1_n8047_22344# m1_n8283_19850# m1_n8283_19850# pfet$29
Xpfet$1_0 vdd vdd m1_3049_25662# m1_2912_25858# pfet$1
Xpfet$1_92 vdd vdd m1_28492_25858# m1_29607_24346# pfet$1
Xpfet$1_81 vdd vdd m1_18339_24542# m1_15943_25858# pfet$1
Xpfet$1_70 vdd vdd m1_14156_24542# m1_11760_25858# pfet$1
Xnfet$14_7 m1_488_21786# m1_488_21786# vss vss m1_n674_21586# vss nfet$14
Xnfet$21_8 m1_3015_15778# m1_3015_15778# m1_2905_18030# m1_2905_18030# m1_3141_17358#
+ vss nfet$21
Xpfet$27_0 vdd vdd m1_n10796_25662# m1_n10933_25858# pfet$27
Xnfet$6_3 m1_9288_21786# vss m1_9418_21590# vss nfet$6
Xpfet$13_6 vdd m1_34278_25658# m1_35071_24542# m1_32330_25662# pfet$13
Xpfet$20_7 vdd m1_27292_16202# m1_26807_17518# m1_27190_17836# pfet$20
Xnfet$4_0 m1_n3534_17714# m1_n3534_17714# vss vss m1_3454_20470# vss nfet$4
Xnfet$14_17 m1_29256_21786# m1_29256_21786# vss vss m1_28094_21586# vss nfet$14
Xnfet$5_75 sd3 vss m1_17697_15478# vss nfet$5
Xnfet$5_64 m1_13668_17714# vss m1_13198_17714# vss nfet$5
Xnfet$5_53 m1_22848_17343# vss m1_23007_17836# vss nfet$5
Xnfet$5_31 m1_1933_17343# m1_3989_15778# m1_3372_16080# vss nfet$5
Xnfet$5_20 m1_1119_17714# vss m1_1709_17518# vss nfet$5
Xnfet$5_42 m1_n811_16080# vss m1_n1168_15778# vss nfet$5
Xnfet$10_1 m1_n789_25858# vss m1_n647_25662# vss nfet$10
Xpfet$3_27 vdd m1_14422_22513# m1_14422_22513# m1_14022_22402# m1_14556_21786# m1_14556_21786#
+ pfet$3
Xpfet$3_16 vdd m1_24973_22513# m1_24973_22513# m1_23945_22102# m1_25739_21786# m1_25739_21786#
+ pfet$3
Xpfet$27_13 vdd vdd m1_n8055_24542# m1_n8625_26174# pfet$27
Xpfet$5_7 vdd vdd m1_4637_21786# m1_4005_21786# pfet$5
Xpfet$1_105 vdd vdd m1_30888_24542# m1_28492_25858# pfet$1
Xnfet$2_76 m1_28492_25858# vss m1_28634_25662# vss nfet$2
Xnfet$2_65 m1_28492_25858# vss m1_25107_21786# vss nfet$2
Xnfet$2_54 m1_24309_25858# vss m1_24451_25662# vss nfet$2
Xnfet$2_43 m1_15461_25858# vss m1_15598_25662# vss nfet$2
Xnfet$2_32 m1_15461_25858# m1_17546_25658# m1_18339_24542# vss nfet$2
Xnfet$2_21 m1_11278_25858# m1_11902_25662# m1_11639_23922# vss nfet$2
Xnfet$2_10 m1_7577_25858# vss m1_9973_24542# vss nfet$2
Xpfet$3_4 vdd vdd vdd m1_9877_22102# m1_9418_21590# m1_9418_21590# pfet$3
Xnfet$22_17 m1_21880_15478# m1_21880_15478# m1_n3206_20274# m1_n3206_20274# m1_23924_20470#
+ vss nfet$22
Xpfet$1_1 vdd m1_3536_25662# m1_3273_23922# m1_3049_25662# pfet$1
Xnfet$28_2 m1_n3206_20274# m1_n3206_20274# vss vss m1_n3724_20470# vss nfet$28
Xnfet$14_8 m1_25739_21786# m1_25739_21786# vss vss m1_24577_21586# vss nfet$14
Xnfet$21_9 m1_2194_16202# m1_2194_16202# vss vss m1_1676_16398# vss nfet$21
Xpfet$27_1 vdd vdd m1_n10309_25662# m1_n10452_25858# pfet$27
Xpfet$1_93 vdd m1_28991_24224# m1_30095_25658# m1_28010_25858# pfet$1
Xpfet$1_82 vdd vdd m1_21241_24346# m1_n7513_20152# pfet$1
Xpfet$1_71 vdd vdd m1_11039_21786# m1_11760_25858# pfet$1
Xpfet$1_60 vdd vdd m1_20126_25858# m1_21241_24346# pfet$1
Xnfet$33_0 m1_n8283_20611# vss m1_n8283_19850# vss nfet$33
Xnfet$6_4 m1_7522_21786# vss m1_8154_21786# vss nfet$6
Xpfet$13_7 vdd m1_32554_23922# m1_32818_24542# m1_32193_25858# pfet$13
Xnfet$4_1 m1_2384_19550# m1_2384_19550# vss vss m1_2822_20470# vss nfet$4
Xnfet$5_76 m1_14482_17343# m1_16538_15778# m1_15921_16080# vss nfet$5
Xnfet$5_65 m1_14482_17343# m1_14743_16202# m1_14258_17518# vss nfet$5
Xnfet$5_54 m1_22848_17343# m1_23109_16202# m1_22624_17518# vss nfet$5
Xnfet$5_32 m1_2092_17836# m1_3015_15778# m1_2194_16202# vss nfet$5
Xnfet$5_21 m1_1933_17343# m1_2194_16202# m1_1709_17518# vss nfet$5
Xnfet$5_10 m1_11738_16080# vss m1_11381_15778# vss nfet$5
Xnfet$5_43 sd8 vss m1_n3218_15478# vss nfet$5
Xnfet$10_2 m1_n1271_25858# vss m1_n1134_25662# vss nfet$10
Xpfet$3_28 vdd m1_14422_22513# m1_14422_22513# m1_13394_22102# m1_15188_21786# m1_15188_21786#
+ pfet$3
Xpfet$3_17 vdd m1_21456_22513# m1_21456_22513# m1_21056_22402# m1_21590_21786# m1_21590_21786#
+ pfet$3
Xpfet$5_8 vdd vdd m1_2384_21590# m1_2254_21786# pfet$5
Xpfet$1_106 vdd vdd m1_25107_21786# m1_28492_25858# pfet$1
Xnfet$2_44 m1_15822_23922# vss m1_16442_24224# vss nfet$2
Xnfet$2_33 m1_11760_25858# vss m1_14156_24542# vss nfet$2
Xnfet$2_22 m1_11760_25858# vss m1_11902_25662# vss nfet$2
Xnfet$2_11 m1_7522_21786# vss m1_11278_25858# vss nfet$2
Xnfet$2_77 m1_28010_25858# vss m1_28147_25662# vss nfet$2
Xnfet$2_66 m1_28010_25858# m1_30095_25658# m1_30888_24542# vss nfet$2
Xnfet$2_55 m1_23827_25858# vss m1_23964_25662# vss nfet$2
Xpfet$3_5 vdd m1_9645_21447# m1_9645_21447# m1_9877_22102# m1_11671_21786# m1_11671_21786#
+ pfet$3
Xnfet$28_3 m1_n6973_21481# m1_n6973_21481# m1_n6839_20152# m1_n6839_20152# m1_n6282_20470#
+ vss nfet$28
Xpfet$1_2 vdd vdd m1_3394_25858# m1_4509_24346# pfet$1
Xnfet$14_9 m1_25107_21786# m1_25107_21786# vss vss m1_23945_21586# vss nfet$14
Xpfet$1_94 vdd m1_28492_25858# vdd m1_30095_25658# pfet$1
Xpfet$1_83 vdd m1_21729_25658# m1_22522_24542# m1_19781_25662# pfet$1
Xpfet$1_72 vdd m1_13363_25658# m1_14156_24542# m1_11415_25662# pfet$1
Xpfet$1_61 vdd m1_24452_24542# vdd m1_25424_24346# pfet$1
Xpfet$1_50 vdd vdd m1_20268_25662# m1_20126_25858# pfet$1
Xnfet$33_1 m1_n7513_20152# m1_n8283_19850# vss vss nfet$33
Xnfet$26_0 m1_n10452_25858# m1_n10452_25858# m1_n7186_25858# m1_n7186_25858# m1_n6629_25502#
+ vss nfet$26
Xpfet$27_2 vdd vdd m1_n9952_24224# m1_n10572_23922# pfet$27
Xnfet$6_5 m1_488_21786# vss m1_1120_21786# vss nfet$6
Xpfet$32_0 vdd vdd vdd m1_n5019_19550# m1_n4485_20152# m1_n4485_20152# pfet$32
Xnfet$4_2 m1_5901_19550# m1_5901_19550# vss vss m1_6339_20470# vss nfet$4
Xnfet$5_77 sd4 vss m1_13514_15478# vss nfet$5
Xnfet$5_66 m1_n7513_20152# vss m1_14127_16080# vss nfet$5
Xnfet$5_55 m1_22034_17714# vss m1_24904_15778# vss nfet$5
Xnfet$5_44 m1_n2091_17836# m1_n811_16080# m1_n1278_18030# vss nfet$5
Xnfet$5_33 sd7 vss m1_965_15478# vss nfet$5
Xnfet$5_22 m1_6116_17343# m1_6377_16202# m1_5892_17518# vss nfet$5
Xnfet$5_11 m1_10299_17343# m1_12355_15778# m1_11738_16080# vss nfet$5
Xnfet$10_3 m1_n7513_20152# vss m1_326_24346# vss nfet$10
Xpfet$3_29 vdd vdd vdd m1_14022_22402# m1_12805_21786# m1_12805_21786# pfet$3
Xpfet$5_9 vdd vdd m1_22222_21786# m1_21590_21786# pfet$5
Xpfet$3_18 vdd vdd vdd m1_24573_22402# m1_23356_21786# m1_23356_21786# pfet$3
Xpfet$1_107 vdd m1_24309_25858# vdd m1_25912_25658# pfet$1
Xnfet$2_78 m1_28010_25858# m1_28634_25662# m1_28371_23922# vss nfet$2
Xnfet$2_67 m1_28492_25858# vss m1_30888_24542# vss nfet$2
Xnfet$2_56 m1_19781_25662# m1_20625_24224# m1_21729_25658# vss nfet$2
Xnfet$2_45 m1_15461_25858# m1_16085_25662# m1_15822_23922# vss nfet$2
Xnfet$2_34 m1_11278_25858# m1_13363_25658# m1_14156_24542# vss nfet$2
Xnfet$2_23 m1_11278_25858# vss m1_11415_25662# vss nfet$2
Xnfet$2_12 m1_7577_25858# vss m1_7522_21786# vss nfet$2
Xpfet$3_6 vdd vdd vdd m1_10505_22402# m1_9288_21786# m1_9288_21786# pfet$3
Xnfet$28_4 m1_2590_19404# m1_2590_19404# vss vss m1_n2445_21430# vss nfet$28
Xpfet$1_3 vdd m1_3394_25858# vdd m1_4997_25658# pfet$1
Xpfet$1_95 vdd vdd m1_28991_24224# m1_28371_23922# pfet$1
Xnfet$19_0 m1_34093_22102# vss fout vss nfet$19
Xpfet$1_84 vdd vdd m1_23827_25858# m1_18073_21786# pfet$1
Xpfet$1_73 vdd m1_16086_24542# vdd m1_17058_24346# pfet$1
Xpfet$1_62 vdd vdd m1_24452_24542# m1_24808_24224# pfet$1
Xpfet$1_51 vdd vdd m1_20625_24224# m1_20005_23922# pfet$1
Xpfet$1_40 vdd vdd m1_11760_25858# m1_12875_24346# pfet$1
Xnfet$33_2 m1_n8145_21908# vss m1_n8283_20611# vss nfet$33
Xpfet$27_3 vdd vdd m1_n4978_24224# vss pfet$27
Xnfet$26_1 m1_n6111_25858# m1_n6111_25858# vss vss m1_n6629_25502# vss nfet$26
Xnfet$6_6 m1_5771_21786# vss m1_5901_21590# vss nfet$6
Xpfet$25_0 vdd vdd m1_n8625_26174# m1_n9336_24346# pfet$25
Xnfet$4_3 m1_4832_17714# m1_4832_17714# vss vss m1_10488_20470# vss nfet$4
Xnfet$5_78 m1_14641_17836# m1_15564_15778# m1_14743_16202# vss nfet$5
Xnfet$5_67 m1_17381_17714# vss m1_14482_17343# vss nfet$5
Xnfet$5_56 m1_24287_16080# vss m1_23930_15778# vss nfet$5
Xnfet$5_45 m1_n3064_17714# vss m1_n194_15778# vss nfet$5
Xnfet$5_34 m1_n2250_17343# vss m1_n2091_17836# vss nfet$5
Xnfet$5_23 m1_5302_17714# vss m1_4832_17714# vss nfet$5
Xnfet$5_12 m1_9485_17714# vss m1_12355_15778# vss nfet$5
Xnfet$10_4 m1_n789_25858# vss m1_1607_24542# vss nfet$10
Xpfet$3_19 vdd m1_24973_22513# m1_24973_22513# m1_24573_22402# m1_25107_21786# m1_25107_21786#
+ pfet$3
Xnfet$2_0 m1_3394_25858# vss m1_5790_24542# vss nfet$2
Xpfet$1_108 vdd vdd m1_25424_24346# m1_n7513_20152# pfet$1
Xnfet$2_79 pd7 vss m1_19839_21786# vss nfet$2
Xnfet$2_68 m1_n7513_20152# vss m1_29607_24346# vss nfet$2
Xnfet$2_57 m1_20126_25858# vss m1_20268_25662# vss nfet$2
Xnfet$2_46 m1_20126_25858# vss m1_18073_21786# vss nfet$2
Xnfet$2_35 m1_15598_25662# m1_15822_23922# m1_16086_24542# vss nfet$2
Xnfet$2_24 m1_7095_25858# m1_7719_25662# m1_7456_23922# vss nfet$2
Xnfet$2_13 m1_11415_25662# m1_11639_23922# m1_11903_24542# vss nfet$2
Xpfet$3_7 vdd m1_354_22513# m1_354_22513# m1_n674_22102# m1_1120_21786# m1_1120_21786#
+ pfet$3
Xpfet$1_4 vdd vdd m1_3893_24224# m1_3273_23922# pfet$1
Xnfet$28_5 m1_6107_19404# m1_6107_19404# m1_n5227_21418# m1_n5227_21418# m1_n2445_21430#
+ vss nfet$28
Xpfet$1_96 vdd m1_28635_24542# vdd m1_29607_24346# pfet$1
Xpfet$1_85 vdd m1_24188_23922# m1_24452_24542# m1_23827_25858# pfet$1
Xpfet$1_74 vdd vdd m1_14556_21786# m1_15943_25858# pfet$1
Xpfet$1_63 vdd vdd m1_19781_25662# m1_19644_25858# pfet$1
Xpfet$1_52 vdd m1_20268_25662# m1_20005_23922# m1_19781_25662# pfet$1
Xpfet$1_41 vdd vdd m1_9288_21786# pd4 pfet$1
Xpfet$1_30 vdd vdd m1_2912_25858# m1_488_21786# pfet$1
Xnfet$33_3 m1_n8283_19850# m1_n8283_20611# vss vss nfet$33
Xpfet$27_4 vdd vdd m1_n5571_25662# m1_n10452_25858# pfet$27
Xnfet$6_7 m1_4005_21786# vss m1_4637_21786# vss nfet$6
Xpfet$18_0 vdd m1_32818_20470# m1_32818_20470# m1_33050_19550# m1_30256_19792# m1_30256_19792#
+ pfet$18
Xnfet$4_4 m1_9418_19550# m1_9418_19550# vss vss m1_9856_20470# vss nfet$4
Xnfet$31_0 m1_n10933_25858# m1_n8848_25658# m1_n8055_24542# vss nfet$31
Xpfet$25_1 vdd m1_n8625_26174# vdd m1_n8848_25658# pfet$25
Xnfet$5_79 m1_15921_16080# vss m1_15564_15778# vss nfet$5
Xnfet$5_68 m1_18665_17343# m1_18926_16202# m1_18441_17518# vss nfet$5
Xnfet$5_57 m1_22848_17343# m1_24904_15778# m1_24287_16080# vss nfet$5
Xnfet$5_46 m1_22034_17714# vss m1_21564_17714# vss nfet$5
Xnfet$5_24 m1_4832_17714# vss m1_1933_17343# vss nfet$5
Xnfet$5_13 m1_10458_17836# m1_11381_15778# m1_10560_16202# vss nfet$5
Xnfet$5_35 m1_n7513_20152# vss m1_5761_16080# vss nfet$5
Xnfet$10_5 m1_n789_25858# vss m1_488_21786# vss nfet$10
Xnfet$2_1 m1_2912_25858# m1_4997_25658# m1_5790_24542# vss nfet$2
Xpfet$1_109 vdd m1_12259_24224# m1_13363_25658# m1_11278_25858# pfet$1
Xnfet$2_69 m1_24309_25858# vss m1_26705_24542# vss nfet$2
Xnfet$2_58 m1_20005_23922# vss m1_20625_24224# vss nfet$2
Xnfet$2_47 m1_23964_25662# m1_24188_23922# m1_24452_24542# vss nfet$2
Xnfet$2_36 m1_11760_25858# vss m1_11039_21786# vss nfet$2
Xnfet$2_25 m1_7232_25662# m1_8076_24224# m1_9180_25658# vss nfet$2
Xnfet$2_14 m1_n7513_20152# vss m1_8692_24346# vss nfet$2
Xpfet$3_8 vdd vdd vdd m1_6360_22102# m1_5901_21590# m1_5901_21590# pfet$3
Xpfet$4_30 vdd vdd vdd m1_24560_19550# m1_21880_15478# m1_21880_15478# pfet$4
Xpfet$1_5 vdd m1_3893_24224# m1_4997_25658# m1_2912_25858# pfet$1
Xnfet$28_6 m1_n5764_21786# m1_n5764_21786# vss vss m1_n6282_21430# vss nfet$28
Xpfet$1_97 vdd vdd m1_21590_21786# m1_24309_25858# pfet$1
Xpfet$1_86 vdd m1_28634_25662# m1_28371_23922# m1_28147_25662# pfet$1
Xpfet$1_75 vdd vdd m1_19644_25858# m1_14556_21786# pfet$1
Xpfet$1_64 vdd vdd m1_22522_24542# m1_20126_25858# pfet$1
Xpfet$1_53 vdd m1_20625_24224# m1_21729_25658# m1_19644_25858# pfet$1
Xpfet$1_42 vdd m1_11760_25858# vdd m1_13363_25658# pfet$1
Xpfet$1_31 vdd m1_3273_23922# m1_3537_24542# m1_2912_25858# pfet$1
Xpfet$1_20 vdd vdd m1_4509_24346# m1_n7513_20152# pfet$1
Xpfet$27_5 vdd vdd m1_n4847_25662# m1_n10452_25858# pfet$27
Xnfet$6_8 m1_2254_21786# vss m1_2384_21590# vss nfet$6
Xpfet$18_1 vdd vdd vdd m1_33050_19550# m1_31535_19792# m1_31535_19792# pfet$18
Xnfet$24_0 m1_n6274_17836# m1_n4994_16080# m1_n5461_18030# vss nfet$24
Xnfet$31_1 m1_n10796_25662# m1_n10572_23922# m1_n10308_24542# vss nfet$31
Xpfet$25_2 vdd m1_n3651_26174# vdd m1_n4978_24224# pfet$25
.ends

.subckt asc_drive_buffer$6 vss in vdd out
Xpfet$69_0 vdd vdd m1_4002_n1060# m1_3466_n454# pfet$69
Xpfet$67_0 out out m1_4274_n1060# vdd m1_4274_n1060# out vdd vdd m1_4274_n1060# out
+ m1_4274_n1060# m1_4274_n1060# out m1_4274_n1060# vdd m1_4274_n1060# vdd m1_4274_n1060#
+ pfet$67
Xnfet$73_0 m1_3466_n454# vss m1_4002_n1060# vss nfet$73
Xnfet$71_0 m1_4274_n1060# vss m1_4002_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ m1_4274_n1060# vss m1_4002_n1060# vss nfet$71
Xpfet$70_0 vdd vdd m1_3466_n454# in pfet$70
Xpfet$68_0 m1_4274_n1060# vdd vdd m1_4274_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ vdd m1_4002_n1060# m1_4002_n1060# pfet$68
Xnfet$74_0 in vss m1_3466_n454# vss nfet$74
Xnfet$72_0 out out vss m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# m1_4274_n1060#
+ m1_4274_n1060# out m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# vss vss
+ nfet$72
.ends

.subckt asc_hysteresis_buffer$10 vss in vdd out
Xnfet$47_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$47
Xnfet$45_0 m1_348_648# vss m1_884_42# vss nfet$45
Xpfet$44_0 vdd vdd m1_884_42# m1_1156_42# pfet$44
Xpfet$42_0 vdd vdd m1_348_648# in pfet$42
Xpfet$40_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd m1_884_42#
+ m1_884_42# pfet$40
Xnfet$48_0 m1_1156_42# vss m1_884_42# vss nfet$48
Xnfet$46_0 in vss m1_348_648# vss nfet$46
Xnfet$44_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$44
Xpfet$43_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$43
Xpfet$41_0 vdd vdd m1_884_42# m1_348_648# pfet$41
.ends

.subckt pfet$37 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$41 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pass1u05u$1 VDD VSS ind ins clkn clkp
Xpfet$37_0 VDD ind ins clkp pfet$37
Xnfet$41_0 clkn ind ins VSS nfet$41
.ends

.subckt nfet$40 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$34 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_954_0# w_n180_n88# a_854_n136#
+ a_n92_0# a_446_n136# a_650_n136# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt pfet$38 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$42 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt inv1u05u$1 in VSS out VDD
Xpfet$38_0 VDD VDD out in pfet$38
Xnfet$42_0 in VSS out VSS nfet$42
.ends

.subckt pfet$36 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=4.55p ps=15.3u w=7u l=0.5u
.ends

.subckt pfet$39 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.5u
.ends

.subckt nfet$38 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt nfet$43 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$35 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_954_0# w_n180_n88#
+ a_38_n60# a_n92_0# a_1058_n60# a_854_n60# a_342_0# a_138_0# a_650_n60#
X0 a_954_0# a_854_n60# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n60# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt nfet$39 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt xp_programmable_basic_pump$1 up vdd s1 s2 s3 s4 down out iref vss
Xpass1u05u$1_2 vdd vss iref pass1u05u$1_2/ins s1 inv1u05u$1_3/out pass1u05u$1
Xnfet$40_6 m1_n7879_n12170# pass1u05u$1_0/ins m1_n7879_n12170# out pass1u05u$1_0/ins
+ vss nfet$40
Xpfet$34_7 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$34
Xpass1u05u$1_3 vdd vss pass1u05u$1_7/ind pass1u05u$1_3/ins s1 inv1u05u$1_3/out pass1u05u$1
Xinv1u05u$1_0 s4 vss inv1u05u$1_0/out vdd inv1u05u$1
Xnfet$40_7 m1_n7879_n12170# pass1u05u$1_0/ins m1_n7879_n12170# out pass1u05u$1_0/ins
+ vss nfet$40
Xpfet$34_8 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$34
Xpass1u05u$1_4 vdd vss pass1u05u$1_7/ind pass1u05u$1_4/ins s2 inv1u05u$1_2/out pass1u05u$1
Xinv1u05u$1_1 s3 vss inv1u05u$1_1/out vdd inv1u05u$1
Xnfet$40_8 vss vdd vss m1_n8144_n9165# vdd vss nfet$40
Xpfet$34_9 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$34
Xpass1u05u$1_5 vdd vss pass1u05u$1_7/ind pass1u05u$1_5/ins s3 inv1u05u$1_1/out pass1u05u$1
Xpfet$36_20 vdd vdd vdd vdd pfet$36
Xpfet$39_0 vdd s3 pass1u05u$1_5/ins vdd pfet$39
Xinv1u05u$1_2 s2 vss inv1u05u$1_2/out vdd inv1u05u$1
Xnfet$40_9 m1_n7216_n8262# iref m1_n7216_n8262# pass1u05u$1_7/ind iref vss nfet$40
Xpass1u05u$1_6 vdd vss iref pass1u05u$1_6/ins s4 inv1u05u$1_0/out pass1u05u$1
Xinv1u05u$1_3 s1 vss inv1u05u$1_3/out vdd inv1u05u$1
Xpfet$36_21 vdd vdd vdd vdd pfet$36
Xpfet$39_1 vdd s2 pass1u05u$1_4/ins vdd pfet$39
Xpass1u05u$1_7 vdd vss pass1u05u$1_7/ind pass1u05u$1_7/ins s4 inv1u05u$1_0/out pass1u05u$1
Xpfet$36_10 vdd vdd vdd vdd pfet$36
Xpfet$39_2 vdd s1 pass1u05u$1_3/ins vdd pfet$39
Xnfet$38_0 pass1u05u$1_6/ins pass1u05u$1_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$38
Xpfet$36_22 vdd vdd vdd vdd pfet$36
Xpfet$36_11 vdd vdd vdd vdd pfet$36
Xpfet$36_23 vdd vdd vdd vdd pfet$36
Xpfet$39_3 vdd s4 pass1u05u$1_7/ins vdd pfet$39
Xnfet$38_1 pass1u05u$1_6/ins pass1u05u$1_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$38
Xpfet$36_12 vdd vdd vdd vdd pfet$36
Xnfet$38_2 pass1u05u$1_6/ins pass1u05u$1_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$38
Xpfet$36_13 vdd vdd vdd vdd pfet$36
Xnfet$43_0 inv1u05u$1_2/out pass1u05u$1_1/ins vss vss nfet$43
Xpfet$36_14 vdd vdd vdd vdd pfet$36
Xnfet$38_3 vss vss vss vss vss vss nfet$38
Xnfet$43_1 inv1u05u$1_3/out pass1u05u$1_2/ins vss vss nfet$43
Xnfet$38_4 pass1u05u$1_6/ins pass1u05u$1_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$38
Xpfet$36_15 vdd vdd vdd vdd pfet$36
Xnfet$43_2 inv1u05u$1_0/out pass1u05u$1_6/ins vss vss nfet$43
Xpfet$35_0 vdd vdd m1_n4127_3649# vss vss m1_n4127_3649# vdd vss vdd vss vss vdd m1_n4127_3649#
+ vss pfet$35
Xpfet$36_16 vdd vdd vdd vdd pfet$36
Xnfet$38_5 vss vss vss vss vss vss nfet$38
Xnfet$43_3 inv1u05u$1_1/out pass1u05u$1_0/ins vss vss nfet$43
Xpfet$35_1 m1_n5580_883# m1_n5580_883# out pass1u05u$1_5/ins pass1u05u$1_5/ins out
+ vdd pass1u05u$1_5/ins m1_n5580_883# pass1u05u$1_5/ins pass1u05u$1_5/ins m1_n5580_883#
+ out pass1u05u$1_5/ins pfet$35
Xpfet$36_17 vdd vdd vdd vdd pfet$36
Xnfet$38_6 pass1u05u$1_6/ins pass1u05u$1_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$38
Xpfet$35_2 m1_n5580_883# m1_n5580_883# out pass1u05u$1_5/ins pass1u05u$1_5/ins out
+ vdd pass1u05u$1_5/ins m1_n5580_883# pass1u05u$1_5/ins pass1u05u$1_5/ins m1_n5580_883#
+ out pass1u05u$1_5/ins pfet$35
Xpfet$36_18 vdd vdd vdd vdd pfet$36
Xnfet$38_7 pass1u05u$1_6/ins pass1u05u$1_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$38
Xpfet$35_3 m1_n5580_883# m1_n5580_883# out pass1u05u$1_5/ins pass1u05u$1_5/ins out
+ vdd pass1u05u$1_5/ins m1_n5580_883# pass1u05u$1_5/ins pass1u05u$1_5/ins m1_n5580_883#
+ out pass1u05u$1_5/ins pfet$35
Xpfet$36_19 vdd vdd vdd vdd pfet$36
Xnfet$38_8 pass1u05u$1_6/ins pass1u05u$1_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$38
Xpfet$35_4 m1_n5580_883# m1_n5580_883# out pass1u05u$1_5/ins pass1u05u$1_5/ins out
+ vdd pass1u05u$1_5/ins m1_n5580_883# pass1u05u$1_5/ins pass1u05u$1_5/ins m1_n5580_883#
+ out pass1u05u$1_5/ins pfet$35
Xnfet$40_10 m1_n8607_n8040# pass1u05u$1_1/ins m1_n8607_n8040# out pass1u05u$1_1/ins
+ vss nfet$40
Xnfet$38_9 pass1u05u$1_6/ins pass1u05u$1_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$38
Xpfet$35_5 m1_n4127_3649# m1_n4127_3649# pass1u05u$1_7/ind pass1u05u$1_7/ind pass1u05u$1_7/ind
+ pass1u05u$1_7/ind vdd pass1u05u$1_7/ind m1_n4127_3649# pass1u05u$1_7/ind pass1u05u$1_7/ind
+ m1_n4127_3649# pass1u05u$1_7/ind pass1u05u$1_7/ind pfet$35
Xnfet$38_10 pass1u05u$1_2/ins pass1u05u$1_2/ins m1_n7679_n8960# m1_n7679_n8960# out
+ vss nfet$38
Xnfet$40_11 m1_n8144_n9165# iref m1_n8144_n9165# iref iref vss nfet$40
Xpfet$34_20 m1_n8156_628# m1_n8156_628# pass1u05u$1_7/ins out out vdd pass1u05u$1_7/ins
+ m1_n8156_628# pass1u05u$1_7/ins pass1u05u$1_7/ins m1_n8156_628# out pass1u05u$1_7/ins
+ pass1u05u$1_7/ins pfet$34
Xnfet$38_11 vss vss vss vss vss vss nfet$38
Xnfet$40_12 vss down vss m1_n8607_n8040# down vss nfet$40
Xpfet$34_21 m1_n6703_2564# m1_n6703_2564# pass1u05u$1_4/ins out out vdd pass1u05u$1_4/ins
+ m1_n6703_2564# pass1u05u$1_4/ins pass1u05u$1_4/ins m1_n6703_2564# out pass1u05u$1_4/ins
+ pass1u05u$1_4/ins pfet$34
Xpfet$34_10 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$34
Xnfet$38_12 down down vss vss m1_n7679_n8960# vss nfet$38
Xnfet$40_13 vss vdd vss m1_n7216_n8262# vdd vss nfet$40
Xpfet$34_22 m1_n8156_628# m1_n8156_628# pass1u05u$1_7/ins out out vdd pass1u05u$1_7/ins
+ m1_n8156_628# pass1u05u$1_7/ins pass1u05u$1_7/ins m1_n8156_628# out pass1u05u$1_7/ins
+ pass1u05u$1_7/ins pfet$34
Xpfet$34_11 vdd vdd up m1_n5450_4559# m1_n5450_4559# vdd up vdd up up vdd m1_n5450_4559#
+ up up pfet$34
Xnfet$38_13 vss vss vss vss vss vss nfet$38
Xnfet$40_14 m1_n8607_n8040# pass1u05u$1_1/ins m1_n8607_n8040# out pass1u05u$1_1/ins
+ vss nfet$40
Xpfet$34_23 m1_n8156_628# m1_n8156_628# pass1u05u$1_7/ins out out vdd pass1u05u$1_7/ins
+ m1_n8156_628# pass1u05u$1_7/ins pass1u05u$1_7/ins m1_n8156_628# out pass1u05u$1_7/ins
+ pass1u05u$1_7/ins pfet$34
Xpfet$34_12 vdd vdd up m1_n6703_2564# m1_n6703_2564# vdd up vdd up up vdd m1_n6703_2564#
+ up up pfet$34
Xnfet$38_14 vss vss vss vss vss vss nfet$38
Xnfet$40_15 vss down vss m1_n8607_n8040# down vss nfet$40
Xpfet$34_24 m1_n5450_4559# m1_n5450_4559# pass1u05u$1_3/ins out out vdd pass1u05u$1_3/ins
+ m1_n5450_4559# pass1u05u$1_3/ins pass1u05u$1_3/ins m1_n5450_4559# out pass1u05u$1_3/ins
+ pass1u05u$1_3/ins pfet$34
Xpfet$34_13 vdd vdd up m1_n6703_2564# m1_n6703_2564# vdd up vdd up up vdd m1_n6703_2564#
+ up up pfet$34
Xnfet$38_15 vss vss vss vss vss vss nfet$38
Xpfet$34_25 m1_n6703_2564# m1_n6703_2564# pass1u05u$1_4/ins out out vdd pass1u05u$1_4/ins
+ m1_n6703_2564# pass1u05u$1_4/ins pass1u05u$1_4/ins m1_n6703_2564# out pass1u05u$1_4/ins
+ pass1u05u$1_4/ins pfet$34
Xpfet$34_14 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$34
Xpfet$34_15 m1_n8156_628# m1_n8156_628# pass1u05u$1_7/ins out out vdd pass1u05u$1_7/ins
+ m1_n8156_628# pass1u05u$1_7/ins pass1u05u$1_7/ins m1_n8156_628# out pass1u05u$1_7/ins
+ pass1u05u$1_7/ins pfet$34
Xnfet$39_0 down down vss vss m1_n8807_n11192# vss nfet$39
Xpfet$34_16 m1_n8156_628# m1_n8156_628# pass1u05u$1_7/ins out out vdd pass1u05u$1_7/ins
+ m1_n8156_628# pass1u05u$1_7/ins pass1u05u$1_7/ins m1_n8156_628# out pass1u05u$1_7/ins
+ pass1u05u$1_7/ins pfet$34
Xnfet$39_1 down down vss vss m1_n8807_n11192# vss nfet$39
Xpfet$34_17 m1_n8156_628# m1_n8156_628# pass1u05u$1_7/ins out out vdd pass1u05u$1_7/ins
+ m1_n8156_628# pass1u05u$1_7/ins pass1u05u$1_7/ins m1_n8156_628# out pass1u05u$1_7/ins
+ pass1u05u$1_7/ins pfet$34
Xpfet$34_18 m1_n8156_628# m1_n8156_628# pass1u05u$1_7/ins out out vdd pass1u05u$1_7/ins
+ m1_n8156_628# pass1u05u$1_7/ins pass1u05u$1_7/ins m1_n8156_628# out pass1u05u$1_7/ins
+ pass1u05u$1_7/ins pfet$34
Xnfet$39_2 down down vss vss m1_n8807_n11192# vss nfet$39
Xnfet$39_3 down down vss vss m1_n8807_n11192# vss nfet$39
Xpfet$34_19 m1_n8156_628# m1_n8156_628# pass1u05u$1_7/ins out out vdd pass1u05u$1_7/ins
+ m1_n8156_628# pass1u05u$1_7/ins pass1u05u$1_7/ins m1_n8156_628# out pass1u05u$1_7/ins
+ pass1u05u$1_7/ins pfet$34
Xnfet$39_4 vss vss vss vss vss vss nfet$39
Xpfet$36_0 vdd vdd vdd vdd pfet$36
Xnfet$39_5 vss vss vss vss vss vss nfet$39
Xnfet$39_10 vss vss vss vss vss vss nfet$39
Xpfet$36_1 vdd vdd vdd vdd pfet$36
Xnfet$39_6 down down vss vss m1_n8807_n11192# vss nfet$39
Xnfet$39_11 vss vss vss vss vss vss nfet$39
Xpfet$36_2 vdd vdd vdd vdd pfet$36
Xnfet$39_7 down down vss vss m1_n8807_n11192# vss nfet$39
Xnfet$39_12 vss vss vss vss vss vss nfet$39
Xpfet$34_0 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$34
Xpfet$36_3 vdd vdd vdd vdd pfet$36
Xnfet$39_8 down down vss vss m1_n8807_n11192# vss nfet$39
Xnfet$39_13 vss vss vss vss vss vss nfet$39
Xpfet$36_4 vdd vdd vdd vdd pfet$36
Xnfet$40_0 m1_n7879_n12170# pass1u05u$1_0/ins m1_n7879_n12170# out pass1u05u$1_0/ins
+ vss nfet$40
Xpfet$34_1 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$34
Xnfet$39_9 down down vss vss m1_n8807_n11192# vss nfet$39
Xnfet$40_1 m1_n7879_n12170# pass1u05u$1_0/ins m1_n7879_n12170# out pass1u05u$1_0/ins
+ vss nfet$40
Xpfet$34_2 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$34
Xpfet$36_5 vdd vdd vdd vdd pfet$36
Xpfet$36_6 vdd vdd vdd vdd pfet$36
Xnfet$40_2 vss down vss m1_n7879_n12170# down vss nfet$40
Xpfet$34_3 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$34
Xpfet$36_7 vdd vdd vdd vdd pfet$36
Xnfet$40_3 vss down vss m1_n7879_n12170# down vss nfet$40
Xpfet$34_4 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$34
Xpass1u05u$1_0 vdd vss iref pass1u05u$1_0/ins s3 inv1u05u$1_1/out pass1u05u$1
Xpfet$36_8 vdd vdd vdd vdd pfet$36
Xnfet$40_4 vss down vss m1_n7879_n12170# down vss nfet$40
Xpfet$34_5 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$34
Xpass1u05u$1_1 vdd vss iref pass1u05u$1_1/ins s2 inv1u05u$1_2/out pass1u05u$1
Xpfet$36_9 vdd vdd vdd vdd pfet$36
Xnfet$40_5 vss down vss m1_n7879_n12170# down vss nfet$40
Xpfet$34_6 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$34
.ends

.subckt nfet$79 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$78 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$84 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$83 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$77 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$76 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt nfet$82 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$75 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$81 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt pfet$74 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$80 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt pfet$72 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$87 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt pfet$79 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt nfet$85 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$78 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$80 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$77 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$83 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt nfet$76 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$82 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt pfet$75 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$81 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$73 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$71 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$88 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$86 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt asc_PFD_DFF_20250831$1 vss fref down up vdd fdiv
Xnfet$79_1 m1_5464_n5483# vss m1_4978_n5483# vss nfet$79
Xpfet$78_0 vdd m1_n5428_n3533# vdd m1_n5650_n4045# pfet$78
Xnfet$84_0 m1_2556_n10129# m1_2556_n10129# vss vss m1_3015_n10205# vss nfet$84
Xpfet$78_1 vdd vdd m1_n5428_n3533# m1_n4678_n3849# pfet$78
Xnfet$84_1 m1_1452_n8889# m1_1452_n8889# m1_1096_n9089# m1_1096_n9089# m1_1550_n9245#
+ vss nfet$84
Xpfet$83_0 vdd m1_5895_n8089# vdd down pfet$83
Xpfet$78_2 vdd m1_n5428_n5842# vdd m1_n5868_n3849# pfet$78
Xnfet$77_0 m1_2779_n3533# vss up vss nfet$77
Xnfet$84_2 m1_2068_n8889# m1_2068_n8889# vss vss m1_1550_n9245# vss nfet$84
Xpfet$78_3 vdd vdd m1_n5428_n5842# m1_n4678_n5482# pfet$78
Xnfet$77_1 m1_2779_n3533# vss m1_3349_n5165# vss nfet$77
Xpfet$83_1 vdd vdd m1_5895_n8089# up pfet$83
Xpfet$76_0 m1_n1926_n4095# vdd vdd m1_n3099_n4095# pfet$76
Xnfet$77_2 m1_2758_n8889# vss m1_2068_n5361# vss nfet$77
Xnfet$84_3 m1_2068_n8889# m1_2068_n8889# m1_2779_n10883# m1_2779_n10883# m1_3015_n10205#
+ vss nfet$84
Xpfet$76_1 m1_n4678_n3849# vdd vdd m1_n1926_n5680# pfet$76
Xnfet$82_0 m1_n4678_n3849# m1_n4678_n3849# m1_n5428_n3533# m1_n5428_n3533# m1_n5192_n4205#
+ vss nfet$82
Xnfet$77_3 m1_832_n5785# vss m1_1452_n5483# vss nfet$77
Xnfet$84_4 m1_n4677_n10522# m1_n4677_n10522# m1_n5427_n10882# m1_n5427_n10882# m1_n5191_n10204#
+ vss nfet$84
Xnfet$75_0 m1_n3885_n4045# m1_832_n5785# m1_1096_n5165# vss nfet$75
Xpfet$76_2 m1_n1926_n5680# vdd vdd m1_n3099_n5680# pfet$76
Xnfet$82_1 m1_n5650_n4045# m1_n5650_n4045# vss vss m1_n5192_n4205# vss nfet$82
Xpfet$81_0 vdd vdd m1_n3098_n10720# m1_n3884_n11124# pfet$81
Xnfet$77_4 vdd vss m1_1095_n4045# vss nfet$77
Xnfet$84_5 m1_n5649_n11124# m1_n5649_n11124# vss vss m1_n5191_n10204# vss nfet$84
Xnfet$75_1 m1_n3885_n4045# m1_1452_n5483# m1_2556_n4049# vss nfet$75
Xpfet$81_1 vdd vdd m1_n3098_n9135# m1_n3884_n9085# pfet$81
Xnfet$82_2 m1_n4678_n5482# m1_n4678_n5482# m1_n5428_n5842# m1_n5428_n5842# m1_n5192_n5164#
+ vss nfet$82
Xpfet$76_3 m1_n4678_n5482# vdd vdd m1_n1926_n4095# pfet$76
Xpfet$74_0 vdd vdd m1_2758_n8889# m1_4978_n5483# pfet$74
Xnfet$84_6 m1_n4677_n8889# m1_n4677_n8889# m1_n5427_n8573# m1_n5427_n8573# m1_n5191_n9245#
+ vss nfet$84
Xnfet$75_2 m1_n3885_n6084# m1_1095_n4045# m1_832_n5785# vss nfet$75
Xnfet$82_3 m1_n5868_n3849# m1_n5868_n3849# vss vss m1_n5192_n5164# vss nfet$82
Xnfet$80_0 m1_n1926_n4095# m1_n3099_n4095# vss vss nfet$80
Xnfet$84_7 m1_n5867_n10544# m1_n5867_n10544# vss vss m1_n5191_n9245# vss nfet$84
Xnfet$75_3 m1_n3885_n6084# m1_2556_n4049# m1_3349_n5165# vss nfet$75
Xnfet$80_1 m1_n4678_n3849# m1_n1926_n5680# vss vss nfet$80
Xnfet$80_2 m1_n1926_n5680# m1_n3099_n5680# vss vss nfet$80
Xpfet$72_0 vdd vdd m1_1096_n5165# m1_1452_n5483# pfet$72
Xnfet$80_3 m1_n4678_n5482# m1_n1926_n4095# vss vss nfet$80
Xpfet$72_1 vdd m1_1096_n5165# vdd m1_2068_n5361# pfet$72
Xpfet$72_2 vdd m1_2779_n3533# vdd m1_2556_n4049# pfet$72
Xpfet$72_3 vdd vdd m1_2779_n3533# m1_2068_n5361# pfet$72
Xnfet$87_0 m1_n4677_n8889# m1_n1925_n10720# vss vss nfet$87
Xnfet$87_1 m1_n1925_n10720# m1_n3098_n10720# vss vss nfet$87
Xnfet$87_2 m1_n4677_n10522# m1_n1925_n9135# vss vss nfet$87
Xpfet$79_0 vdd vdd m1_n3099_n4095# m1_n3885_n4045# pfet$79
Xnfet$85_0 m1_n3884_n9085# m1_1095_n11125# m1_832_n8573# vss nfet$85
Xnfet$87_3 m1_n1925_n9135# m1_n3098_n9135# vss vss nfet$87
Xpfet$79_1 vdd vdd m1_n3099_n5680# m1_n3885_n6084# pfet$79
Xnfet$85_1 m1_n3884_n11124# m1_1452_n8889# m1_2556_n10129# vss nfet$85
Xnfet$78_0 m1_4978_n5483# vss m1_2758_n8889# vss nfet$78
Xpfet$80_20 vdd m1_n5427_n8573# vdd m1_n5867_n10544# pfet$80
Xnfet$85_2 m1_832_n8573# vss m1_1452_n8889# vss nfet$85
Xpfet$77_0 vdd vdd m1_n3885_n4045# m1_n5428_n3533# pfet$77
Xpfet$80_10 vdd vdd m1_3349_n9089# m1_2779_n10883# pfet$80
Xnfet$85_3 vdd vss m1_1095_n11125# vss nfet$85
Xnfet$83_0 m1_n3885_n4045# vss m1_n3099_n4095# vss nfet$83
Xpfet$77_1 vdd vdd m1_n5650_n4045# m1_n5868_n3849# pfet$77
Xpfet$80_11 vdd vdd down m1_2779_n10883# pfet$80
Xnfet$76_0 m1_2068_n5361# m1_2068_n5361# vss vss m1_1550_n5165# vss nfet$76
Xnfet$85_4 m1_n3884_n11124# m1_832_n8573# m1_1096_n9089# vss nfet$85
Xnfet$83_1 m1_n3885_n6084# vss m1_n3099_n5680# vss nfet$83
Xpfet$77_2 vdd vdd m1_n3885_n6084# m1_n5428_n5842# pfet$77
Xpfet$82_0 m1_n4677_n8889# vdd vdd m1_n1925_n10720# pfet$82
Xpfet$80_12 vdd m1_2556_n10129# m1_3349_n9089# m1_n3884_n11124# pfet$80
Xnfet$85_5 m1_2758_n8889# vss m1_2068_n8889# vss nfet$85
Xnfet$76_1 m1_1452_n5483# m1_1452_n5483# m1_1096_n5165# m1_1096_n5165# m1_1550_n5165#
+ vss nfet$76
Xpfet$77_3 vdd vdd m1_n5868_n3849# fref pfet$77
Xpfet$82_1 m1_n1925_n10720# vdd vdd m1_n3098_n10720# pfet$82
Xpfet$75_0 vdd vdd m1_5464_n5483# m1_5895_n8089# pfet$75
Xpfet$80_13 vdd vdd m1_n5427_n8573# m1_n4677_n8889# pfet$80
Xnfet$76_2 m1_2556_n4049# m1_2556_n4049# vss vss m1_3015_n4205# vss nfet$76
Xnfet$85_6 m1_2779_n10883# vss down vss nfet$85
Xpfet$82_2 m1_n4677_n10522# vdd vdd m1_n1925_n9135# pfet$82
Xnfet$81_0 m1_n5428_n3533# vss m1_n3885_n4045# vss nfet$81
Xpfet$75_1 vdd vdd m1_4978_n5483# m1_5464_n5483# pfet$75
Xpfet$80_14 vdd vdd m1_n3884_n11124# m1_n5427_n10882# pfet$80
Xnfet$85_7 m1_2779_n10883# vss m1_3349_n9089# vss nfet$85
Xnfet$76_3 m1_2068_n5361# m1_2068_n5361# m1_2779_n3533# m1_2779_n3533# m1_3015_n4205#
+ vss nfet$76
Xpfet$80_0 vdd vdd m1_2779_n10883# m1_2068_n8889# pfet$80
Xpfet$82_3 m1_n1925_n9135# vdd vdd m1_n3098_n9135# pfet$82
Xnfet$81_1 m1_n5868_n3849# vss m1_n5650_n4045# vss nfet$81
Xpfet$80_15 vdd m1_n5427_n10882# vdd m1_n5649_n11124# pfet$80
Xnfet$85_8 m1_n3884_n9085# m1_2556_n10129# m1_3349_n9089# vss nfet$85
Xnfet$81_2 m1_n5428_n5842# vss m1_n3885_n6084# vss nfet$81
Xpfet$80_1 vdd m1_2779_n10883# vdd m1_2556_n10129# pfet$80
Xpfet$80_16 vdd vdd m1_n5427_n10882# m1_n4677_n10522# pfet$80
Xpfet$73_0 vdd vdd m1_3349_n5165# m1_2779_n3533# pfet$73
Xnfet$85_9 m1_n5427_n10882# vss m1_n3884_n11124# vss nfet$85
Xpfet$80_2 vdd m1_1095_n11125# m1_832_n8573# m1_n3884_n11124# pfet$80
Xnfet$81_3 fref vss m1_n5868_n3849# vss nfet$81
Xpfet$73_1 vdd vdd up m1_2779_n3533# pfet$73
Xpfet$80_17 vdd vdd m1_n5649_n11124# m1_n5867_n10544# pfet$80
Xpfet$73_2 vdd vdd m1_2068_n5361# m1_2758_n8889# pfet$73
Xpfet$80_3 vdd m1_1452_n8889# m1_2556_n10129# m1_n3884_n9085# pfet$80
Xpfet$80_18 vdd vdd m1_n5867_n10544# fdiv pfet$80
Xpfet$80_4 vdd vdd m1_1452_n8889# m1_832_n8573# pfet$80
Xpfet$73_3 vdd vdd m1_1452_n5483# m1_832_n5785# pfet$73
Xpfet$71_0 vdd m1_832_n5785# m1_1096_n5165# m1_n3885_n6084# pfet$71
Xpfet$80_19 vdd vdd m1_n3884_n9085# m1_n5427_n8573# pfet$80
Xpfet$73_4 vdd vdd m1_1095_n4045# vdd pfet$73
Xpfet$80_5 vdd vdd m1_1095_n11125# vdd pfet$80
Xpfet$71_1 vdd m1_1452_n5483# m1_2556_n4049# m1_n3885_n6084# pfet$71
Xnfet$88_0 up up m1_5895_n8089# m1_5895_n8089# m1_5043_n9245# vss nfet$88
Xnfet$85_10 m1_n5867_n10544# vss m1_n5649_n11124# vss nfet$85
Xpfet$71_2 vdd m1_1095_n4045# m1_832_n5785# m1_n3885_n4045# pfet$71
Xpfet$80_6 vdd vdd m1_1096_n9089# m1_1452_n8889# pfet$80
Xnfet$88_1 down down vss vss m1_5043_n9245# vss nfet$88
Xnfet$85_11 fdiv vss m1_n5867_n10544# vss nfet$85
Xpfet$80_7 vdd m1_832_n8573# m1_1096_n9089# m1_n3884_n9085# pfet$80
Xpfet$71_3 vdd m1_2556_n4049# m1_3349_n5165# m1_n3885_n4045# pfet$71
Xnfet$85_12 m1_n5427_n8573# vss m1_n3884_n9085# vss nfet$85
Xpfet$80_8 vdd m1_1096_n9089# vdd m1_2068_n8889# pfet$80
Xpfet$80_9 vdd vdd m1_2068_n8889# m1_2758_n8889# pfet$80
Xnfet$86_0 m1_n3884_n11124# vss m1_n3098_n10720# vss nfet$86
Xnfet$86_1 m1_n3884_n9085# vss m1_n3098_n9135# vss nfet$86
Xnfet$79_0 m1_5895_n8089# vss m1_5464_n5483# vss nfet$79
.ends

.subckt nfet$68 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt nfet$66 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$65 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$63 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$69 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$67 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$66 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$64 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$70 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$62 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt asc_drive_buffer_up$1 vss out in vdd
Xnfet$68_0 m1_n30_1318# vss m1_506_712# vss nfet$68
Xnfet$66_0 m1_778_712# vss m1_506_712# m1_506_712# m1_506_712# m1_778_712# m1_778_712#
+ vss m1_506_712# vss nfet$66
Xpfet$65_0 vdd vdd m1_n30_1318# m1_n566_1318# pfet$65
Xpfet$63_0 m1_778_712# vdd vdd m1_778_712# m1_506_712# m1_506_712# m1_778_712# vdd
+ m1_506_712# m1_506_712# pfet$63
Xnfet$69_0 m1_n566_1318# vss m1_n30_1318# vss nfet$69
Xnfet$67_0 out out vss m1_778_712# m1_778_712# out vss m1_778_712# m1_778_712# m1_778_712#
+ out m1_778_712# m1_778_712# out vss m1_778_712# vss vss nfet$67
Xpfet$66_0 vdd vdd m1_n566_1318# in pfet$66
Xpfet$64_0 vdd vdd m1_506_712# m1_n30_1318# pfet$64
Xnfet$70_0 in vss m1_n566_1318# vss nfet$70
Xpfet$62_0 out out m1_778_712# vdd m1_778_712# out vdd vdd m1_778_712# out m1_778_712#
+ m1_778_712# out m1_778_712# vdd m1_778_712# vdd m1_778_712# pfet$62
.ends

.subckt pfet$84 a_254_0# a_348_560# w_n180_n88# a_414_0# a_n92_0# a_94_0# a_574_0#
+ a_508_560# a_188_560# a_28_560#
X0 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$89 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt BIAS$1 vdd vss 100n 200n res 200p1 200p2
Xpfet$84_13 vdd res vdd res vdd res vdd res res res pfet$84
Xpfet$84_15 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$84
Xpfet$84_14 vdd res vdd 200n vdd 200n vdd res res res pfet$84
Xnfet$89_1 vss vss vss vss vss vss vss vss vss vss nfet$89
Xnfet$89_0 m1_27_n1423# vss 200p1 m1_27_n1423# vss 200p1 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$89
Xnfet$89_2 m1_27_n1423# vss 200p2 m1_27_n1423# vss 200p2 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$89
Xnfet$89_3 vss vss vss vss vss vss vss vss vss vss nfet$89
Xnfet$89_4 m1_27_n1423# vss 200p2 m1_27_n1423# vss 200p2 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$89
Xnfet$89_5 m1_27_n1423# vss 200p1 m1_27_n1423# vss 200p1 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$89
Xnfet$89_6 m1_27_n1423# vss m1_27_n1423# m1_27_n1423# vss m1_27_n1423# m1_27_n1423#
+ vss m1_27_n1423# vss nfet$89
Xnfet$89_7 m1_27_n1423# vss m1_27_n1423# m1_27_n1423# vss m1_27_n1423# m1_27_n1423#
+ vss m1_27_n1423# vss nfet$89
Xpfet$84_0 vdd res vdd 200n vdd 200n vdd res res res pfet$84
Xpfet$84_1 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$84
Xpfet$84_2 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$84
Xpfet$84_3 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$84
Xpfet$84_4 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$84
Xpfet$84_5 vdd res vdd 200n vdd 200n vdd res res res pfet$84
Xpfet$84_6 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$84
Xpfet$84_8 vdd res vdd res vdd res vdd res res res pfet$84
Xpfet$84_7 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$84
Xpfet$84_9 vdd res vdd 100n vdd 100n vdd res res res pfet$84
Xpfet$84_10 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$84
Xpfet$84_11 vdd res vdd 200n vdd 200n vdd res res res pfet$84
Xpfet$84_12 vdd res vdd 100n vdd 100n vdd res res res pfet$84
.ends

.subckt nfet$58 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$49 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$56 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$54 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$48 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$55 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$53 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$46 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$52 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$51 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$50 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt nfet$59 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$58 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$57 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$56 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$49 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$62 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$55 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$54 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$47 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$60 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$53 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$52 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$45 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$51 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$50 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$59 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$57 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$63 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$61 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_lock_detector_20250826$1 ref vdd div vss lock
Xnfet$58_6 m1_17926_34# vss m1_19469_1832# vss nfet$58
Xnfet$49_2 m1_12790_n340# m1_12790_n340# vss m1_11642_n340# m1_11642_n340# m1_12790_n340#
+ vss m1_11642_n340# m1_11642_n340# m1_11642_n340# m1_12790_n340# m1_11642_n340# m1_11642_n340#
+ m1_12790_n340# vss m1_11642_n340# vss vss nfet$49
Xnfet$56_3 m1_15755_n208# m1_15979_2344# m1_16243_1828# vss nfet$56
Xnfet$54_0 m1_n7214_4493# vss m1_n7486_4493# m1_n7486_4493# m1_n7486_4493# m1_n7214_4493#
+ m1_n7214_4493# vss m1_n7486_4493# vss nfet$54
Xpfet$48_1 m1_11642_n340# vdd vdd m1_11642_n340# m1_11370_n340# m1_11370_n340# m1_11642_n340#
+ vdd m1_11370_n340# m1_11370_n340# pfet$48
Xpfet$55_2 vdd vdd m1_n12216_5099# m1_n14454_7868# pfet$55
Xnfet$58_7 vss vss m1_17215_5644# vss nfet$58
Xnfet$54_1 m1_n15602_4493# vss m1_n15874_4493# m1_n15874_4493# m1_n15874_4493# m1_n15602_4493#
+ m1_n15602_4493# vss m1_n15874_4493# vss nfet$54
Xnfet$56_4 m1_15618_7156# m1_17703_6956# m1_18496_5840# vss nfet$56
Xpfet$48_2 m1_3254_n340# vdd vdd m1_3254_n340# m1_2982_n340# m1_2982_n340# m1_3254_n340#
+ vdd m1_2982_n340# m1_2982_n340# pfet$48
Xnfet$49_3 m1_208_n340# m1_208_n340# vss m1_n940_n340# m1_n940_n340# m1_208_n340#
+ vss m1_n940_n340# m1_n940_n340# m1_n940_n340# m1_208_n340# m1_n940_n340# m1_n940_n340#
+ m1_208_n340# vss m1_n940_n340# vss vss nfet$49
Xpfet$53_0 m1_n11408_4493# vdd vdd m1_n11408_4493# m1_n11680_4493# m1_n11680_4493#
+ m1_n11408_4493# vdd m1_n11680_4493# m1_n11680_4493# pfet$53
Xnfet$49_4 m1_12790_7868# m1_12790_7868# vss m1_11642_4493# m1_11642_4493# m1_12790_7868#
+ vss m1_11642_4493# m1_11642_4493# m1_11642_4493# m1_12790_7868# m1_11642_4493# m1_11642_4493#
+ m1_12790_7868# vss m1_11642_4493# vss vss nfet$49
Xnfet$56_5 m1_15755_6960# m1_15979_5220# m1_16243_5840# vss nfet$56
Xnfet$58_8 m1_17926_7472# vss m1_19469_4920# vss nfet$58
Xnfet$54_2 m1_n11408_4493# vss m1_n11680_4493# m1_n11680_4493# m1_n11680_4493# m1_n11408_4493#
+ m1_n11408_4493# vss m1_n11680_4493# vss nfet$54
Xpfet$46_0 vdd vdd m1_7176_n340# m1_6640_1478# pfet$46
Xpfet$48_3 m1_n940_n340# vdd vdd m1_n940_n340# m1_n1212_n340# m1_n1212_n340# m1_n940_n340#
+ vdd m1_n1212_n340# m1_n1212_n340# pfet$48
Xpfet$53_1 m1_n7214_4493# vdd vdd m1_n7214_4493# m1_n7486_4493# m1_n7486_4493# m1_n7214_4493#
+ vdd m1_n7486_4493# m1_n7486_4493# pfet$53
Xnfet$58_9 m1_17926_7472# vss m1_18496_5840# vss nfet$58
Xnfet$49_5 m1_8596_7868# m1_8596_7868# vss m1_7448_4493# m1_7448_4493# m1_8596_7868#
+ vss m1_7448_4493# m1_7448_4493# m1_7448_4493# m1_8596_7868# m1_7448_4493# m1_7448_4493#
+ m1_8596_7868# vss m1_7448_4493# vss vss nfet$49
Xnfet$56_6 m1_15618_7156# m1_16242_6960# m1_15979_5220# vss nfet$56
Xpfet$48_4 m1_n940_4493# vdd vdd m1_n940_4493# m1_n1212_4493# m1_n1212_4493# m1_n940_4493#
+ vdd m1_n1212_4493# m1_n1212_4493# pfet$48
Xnfet$52_0 m1_n6066_7868# m1_n6066_7868# vss m1_n7214_4493# m1_n7214_4493# m1_n6066_7868#
+ vss m1_n7214_4493# m1_n7214_4493# m1_n7214_4493# m1_n6066_7868# m1_n7214_4493# m1_n7214_4493#
+ m1_n6066_7868# vss m1_n7214_4493# vss vss nfet$52
Xpfet$46_1 vdd vdd m1_11370_n340# m1_10834_1478# pfet$46
Xpfet$53_2 m1_n15602_4493# vdd vdd m1_n15602_4493# m1_n15874_4493# m1_n15874_4493#
+ m1_n15602_4493# vdd m1_n15874_4493# m1_n15874_4493# pfet$53
Xnfet$49_6 m1_208_7868# m1_208_7868# vss m1_n940_4493# m1_n940_4493# m1_208_7868#
+ vss m1_n940_4493# m1_n940_4493# m1_n940_4493# m1_208_7868# m1_n940_4493# m1_n940_4493#
+ m1_208_7868# vss m1_n940_4493# vss vss nfet$49
Xnfet$56_7 m1_15755_6960# m1_16599_5522# m1_17703_6956# vss nfet$56
Xpfet$48_5 m1_11642_4493# vdd vdd m1_11642_4493# m1_11370_4493# m1_11370_4493# m1_11642_4493#
+ vdd m1_11370_4493# m1_11370_4493# pfet$48
Xnfet$52_1 m1_n14454_7868# m1_n14454_7868# vss m1_n15602_4493# m1_n15602_4493# m1_n14454_7868#
+ vss m1_n15602_4493# m1_n15602_4493# m1_n15602_4493# m1_n14454_7868# m1_n15602_4493#
+ m1_n15602_4493# m1_n14454_7868# vss m1_n15602_4493# vss vss nfet$52
Xpfet$51_0 vdd m1_17926_34# vdd m1_17703_788# pfet$51
Xpfet$46_2 vdd vdd m1_2982_n340# m1_2446_1478# pfet$46
Xnfet$49_7 m1_4402_7868# m1_4402_7868# vss m1_3254_4493# m1_3254_4493# m1_4402_7868#
+ vss m1_3254_4493# m1_3254_4493# m1_3254_4493# m1_4402_7868# m1_3254_4493# m1_3254_4493#
+ m1_4402_7868# vss m1_3254_4493# vss vss nfet$49
Xpfet$48_6 m1_3254_4493# vdd vdd m1_3254_4493# m1_2982_4493# m1_2982_4493# m1_3254_4493#
+ vdd m1_2982_4493# m1_2982_4493# pfet$48
Xnfet$52_2 m1_n10260_7868# m1_n10260_7868# vss m1_n11408_4493# m1_n11408_4493# m1_n10260_7868#
+ vss m1_n11408_4493# m1_n11408_4493# m1_n11408_4493# m1_n10260_7868# m1_n11408_4493#
+ m1_n11408_4493# m1_n10260_7868# vss m1_n11408_4493# vss vss nfet$52
Xpfet$46_3 vdd vdd m1_n1212_n340# m1_n1748_1478# pfet$46
Xpfet$51_1 vdd vdd m1_17926_34# m1_17215_2028# pfet$51
Xpfet$48_7 m1_7448_4493# vdd vdd m1_7448_4493# m1_7176_4493# m1_7176_4493# m1_7448_4493#
+ vdd m1_7176_4493# m1_7176_4493# pfet$48
Xnfet$50_0 m1_10834_1478# vss m1_11370_n340# vss nfet$50
Xpfet$51_2 vdd m1_16243_1828# vdd m1_17215_2028# pfet$51
Xpfet$46_4 vdd vdd m1_n1212_4493# m1_n1748_5099# pfet$46
Xpfet$46_5 vdd vdd m1_2982_4493# m1_2446_5099# pfet$46
Xnfet$50_1 m1_2446_1478# vss m1_2982_n340# vss nfet$50
Xpfet$51_3 vdd vdd m1_16243_1828# m1_16599_2028# pfet$51
Xpfet$46_6 vdd vdd m1_7176_4493# m1_6640_5099# pfet$46
Xnfet$50_2 m1_6640_1478# vss m1_7176_n340# vss nfet$50
Xpfet$51_4 vdd m1_16243_5840# vdd m1_17215_5644# pfet$51
Xpfet$46_7 vdd vdd m1_11370_4493# m1_10834_5099# pfet$46
Xpfet$51_5 vdd vdd m1_16243_5840# m1_16599_5522# pfet$51
Xnfet$50_3 m1_n1748_1478# vss m1_n1212_n340# vss nfet$50
Xnfet$59_0 m1_n14454_7868# vss m1_n12216_5099# vss nfet$59
Xnfet$50_4 m1_10834_5099# vss m1_11370_4493# vss nfet$50
Xpfet$51_6 vdd m1_17926_7472# vdd m1_17703_6956# pfet$51
Xnfet$59_1 div vss m1_n16410_5099# vss nfet$59
Xnfet$50_5 m1_6640_5099# vss m1_7176_4493# vss nfet$50
Xpfet$51_7 vdd vdd m1_17926_7472# m1_17215_5644# pfet$51
Xpfet$58_0 vdd m1_19675_2344# vdd m1_19469_1832# pfet$58
Xpfet$58_1 vdd vdd m1_19675_2344# m1_19469_4920# pfet$58
Xnfet$59_2 m1_n10260_7868# vss m1_n8022_5099# vss nfet$59
Xnfet$50_6 m1_n1748_5099# vss m1_n1212_4493# vss nfet$50
Xnfet$50_7 m1_2446_5099# vss m1_2982_4493# vss nfet$50
Xnfet$57_0 m1_17215_2028# m1_17215_2028# m1_17926_34# m1_17926_34# m1_18162_712# vss
+ nfet$57
Xnfet$57_1 m1_17703_788# m1_17703_788# vss vss m1_18162_712# vss nfet$57
Xpfet$56_0 vdd vdd vdd m1_n3798_6028# div div pfet$56
Xnfet$57_2 m1_16599_2028# m1_16599_2028# m1_16243_1828# m1_16243_1828# m1_16697_1672#
+ vss nfet$57
Xpfet$49_0 vdd vdd m1_16599_2028# m1_15979_2344# pfet$49
Xnfet$62_0 m1_19469_4920# m1_19469_4920# m1_19675_2344# m1_19675_2344# m1_19911_1672#
+ vss nfet$62
Xpfet$56_1 vdd m1_n4030_5270# m1_n4030_5270# m1_n3798_6028# m1_n6066_7868# m1_n6066_7868#
+ pfet$56
Xnfet$57_3 m1_17215_2028# m1_17215_2028# vss vss m1_16697_1672# vss nfet$57
Xpfet$49_1 vdd vdd m1_16242_n208# m1_n2336_5099# pfet$49
Xnfet$55_0 m1_8596_n340# vss m1_10834_1478# vss nfet$55
Xnfet$62_1 m1_19469_1832# m1_19469_1832# vss vss m1_19911_1672# vss nfet$62
Xnfet$57_4 m1_17215_5644# m1_17215_5644# vss vss m1_16697_5840# vss nfet$57
Xpfet$49_2 vdd vdd m1_15755_n208# m1_15618_394# pfet$49
Xnfet$55_1 m1_4402_n340# vss m1_6640_1478# vss nfet$55
Xpfet$54_0 vdd vdd m1_n11680_4493# m1_n12216_5099# pfet$54
Xnfet$57_5 m1_16599_5522# m1_16599_5522# m1_16243_5840# m1_16243_5840# m1_16697_5840#
+ vss nfet$57
Xpfet$49_3 vdd vdd m1_18496_1828# m1_17926_34# pfet$49
Xnfet$55_2 ref vss m1_n1748_1478# vss nfet$55
Xpfet$47_0 m1_8596_n340# m1_8596_n340# m1_7448_n340# vdd m1_7448_n340# m1_8596_n340#
+ vdd vdd m1_7448_n340# m1_8596_n340# m1_7448_n340# m1_7448_n340# m1_8596_n340# m1_7448_n340#
+ vdd m1_7448_n340# vdd m1_7448_n340# pfet$47
Xnfet$60_0 div m1_n4030_5270# vss vss nfet$60
Xpfet$54_1 vdd vdd m1_n7486_4493# m1_n8022_5099# pfet$54
Xnfet$57_6 m1_17215_5644# m1_17215_5644# m1_17926_7472# m1_17926_7472# m1_18162_6800#
+ vss nfet$57
Xnfet$53_0 m1_n8022_5099# vss m1_n7486_4493# vss nfet$53
Xpfet$49_4 vdd vdd m1_15618_394# m1_12790_n340# pfet$49
Xpfet$47_1 m1_12790_n340# m1_12790_n340# m1_11642_n340# vdd m1_11642_n340# m1_12790_n340#
+ vdd vdd m1_11642_n340# m1_12790_n340# m1_11642_n340# m1_11642_n340# m1_12790_n340#
+ m1_11642_n340# vdd m1_11642_n340# vdd m1_11642_n340# pfet$47
Xnfet$60_1 m1_n6066_7868# vss m1_n4030_5270# vss nfet$60
Xnfet$55_3 m1_n2336_5099# vss m1_n1748_5099# vss nfet$55
Xpfet$54_2 vdd vdd m1_n15874_4493# m1_n16410_5099# pfet$54
Xnfet$57_7 m1_17703_6956# m1_17703_6956# vss vss m1_18162_6800# vss nfet$57
Xnfet$55_4 m1_8596_7868# vss m1_10834_5099# vss nfet$55
Xpfet$49_5 vdd vdd m1_17215_2028# vss pfet$49
Xnfet$53_1 m1_n16410_5099# vss m1_n15874_4493# vss nfet$53
Xpfet$47_2 m1_4402_n340# m1_4402_n340# m1_3254_n340# vdd m1_3254_n340# m1_4402_n340#
+ vdd vdd m1_3254_n340# m1_4402_n340# m1_3254_n340# m1_3254_n340# m1_4402_n340# m1_3254_n340#
+ vdd m1_3254_n340# vdd m1_3254_n340# pfet$47
Xpfet$52_0 m1_n10260_7868# m1_n10260_7868# m1_n11408_4493# vdd m1_n11408_4493# m1_n10260_7868#
+ vdd vdd m1_n11408_4493# m1_n10260_7868# m1_n11408_4493# m1_n11408_4493# m1_n10260_7868#
+ m1_n11408_4493# vdd m1_n11408_4493# vdd m1_n11408_4493# pfet$52
Xnfet$55_5 m1_4402_7868# vss m1_6640_5099# vss nfet$55
Xpfet$49_6 vdd vdd m1_19469_1832# m1_17926_34# pfet$49
Xpfet$47_3 m1_208_n340# m1_208_n340# m1_n940_n340# vdd m1_n940_n340# m1_208_n340#
+ vdd vdd m1_n940_n340# m1_208_n340# m1_n940_n340# m1_n940_n340# m1_208_n340# m1_n940_n340#
+ vdd m1_n940_n340# vdd m1_n940_n340# pfet$47
Xnfet$53_2 m1_n12216_5099# vss m1_n11680_4493# vss nfet$53
Xpfet$45_0 vdd vdd m1_6640_1478# m1_4402_n340# pfet$45
Xpfet$52_1 m1_n6066_7868# m1_n6066_7868# m1_n7214_4493# vdd m1_n7214_4493# m1_n6066_7868#
+ vdd vdd m1_n7214_4493# m1_n6066_7868# m1_n7214_4493# m1_n7214_4493# m1_n6066_7868#
+ m1_n7214_4493# vdd m1_n7214_4493# vdd m1_n7214_4493# pfet$52
Xnfet$55_6 m1_208_n340# vss m1_2446_1478# vss nfet$55
Xpfet$49_7 vdd vdd m1_17215_5644# vss pfet$49
Xpfet$47_4 m1_208_7868# m1_208_7868# m1_n940_4493# vdd m1_n940_4493# m1_208_7868#
+ vdd vdd m1_n940_4493# m1_208_7868# m1_n940_4493# m1_n940_4493# m1_208_7868# m1_n940_4493#
+ vdd m1_n940_4493# vdd m1_n940_4493# pfet$47
Xnfet$51_0 m1_3254_n340# vss m1_2982_n340# m1_2982_n340# m1_2982_n340# m1_3254_n340#
+ m1_3254_n340# vss m1_2982_n340# vss nfet$51
Xpfet$45_1 vdd vdd m1_10834_1478# m1_8596_n340# pfet$45
Xpfet$52_2 m1_n14454_7868# m1_n14454_7868# m1_n15602_4493# vdd m1_n15602_4493# m1_n14454_7868#
+ vdd vdd m1_n15602_4493# m1_n14454_7868# m1_n15602_4493# m1_n15602_4493# m1_n14454_7868#
+ m1_n15602_4493# vdd m1_n15602_4493# vdd m1_n15602_4493# pfet$52
Xnfet$55_7 m1_208_7868# vss m1_2446_5099# vss nfet$55
Xpfet$49_8 vdd vdd m1_19469_4920# m1_17926_7472# pfet$49
Xpfet$47_5 m1_12790_7868# m1_12790_7868# m1_11642_4493# vdd m1_11642_4493# m1_12790_7868#
+ vdd vdd m1_11642_4493# m1_12790_7868# m1_11642_4493# m1_11642_4493# m1_12790_7868#
+ m1_11642_4493# vdd m1_11642_4493# vdd m1_11642_4493# pfet$47
Xnfet$51_1 m1_7448_n340# vss m1_7176_n340# m1_7176_n340# m1_7176_n340# m1_7448_n340#
+ m1_7448_n340# vss m1_7176_n340# vss nfet$51
Xpfet$45_2 vdd vdd m1_n1748_1478# ref pfet$45
Xpfet$50_0 vdd m1_16599_2028# m1_17703_788# m1_15618_394# pfet$50
Xpfet$49_9 vdd vdd m1_18496_5840# m1_17926_7472# pfet$49
Xpfet$47_6 m1_4402_7868# m1_4402_7868# m1_3254_4493# vdd m1_3254_4493# m1_4402_7868#
+ vdd vdd m1_3254_4493# m1_4402_7868# m1_3254_4493# m1_3254_4493# m1_4402_7868# m1_3254_4493#
+ vdd m1_3254_4493# vdd m1_3254_4493# pfet$47
Xpfet$50_1 vdd m1_16242_n208# m1_15979_2344# m1_15755_n208# pfet$50
Xnfet$51_2 m1_11642_n340# vss m1_11370_n340# m1_11370_n340# m1_11370_n340# m1_11642_n340#
+ m1_11642_n340# vss m1_11370_n340# vss nfet$51
Xpfet$45_3 vdd vdd m1_n1748_5099# m1_n2336_5099# pfet$45
Xpfet$47_7 m1_8596_7868# m1_8596_7868# m1_7448_4493# vdd m1_7448_4493# m1_8596_7868#
+ vdd vdd m1_7448_4493# m1_8596_7868# m1_7448_4493# m1_7448_4493# m1_8596_7868# m1_7448_4493#
+ vdd m1_7448_4493# vdd m1_7448_4493# pfet$47
Xpfet$45_4 vdd vdd m1_6640_5099# m1_4402_7868# pfet$45
Xnfet$51_3 m1_n940_n340# vss m1_n1212_n340# m1_n1212_n340# m1_n1212_n340# m1_n940_n340#
+ m1_n940_n340# vss m1_n1212_n340# vss nfet$51
Xpfet$50_2 vdd m1_15979_2344# m1_16243_1828# m1_15618_394# pfet$50
Xnfet$51_4 m1_11642_4493# vss m1_11370_4493# m1_11370_4493# m1_11370_4493# m1_11642_4493#
+ m1_11642_4493# vss m1_11370_4493# vss nfet$51
Xpfet$45_5 vdd vdd m1_10834_5099# m1_8596_7868# pfet$45
Xpfet$50_3 vdd m1_17703_788# m1_18496_1828# m1_15755_n208# pfet$50
Xpfet$45_6 vdd vdd m1_2446_5099# m1_208_7868# pfet$45
Xnfet$51_5 m1_7448_4493# vss m1_7176_4493# m1_7176_4493# m1_7176_4493# m1_7448_4493#
+ m1_7448_4493# vss m1_7176_4493# vss nfet$51
Xpfet$59_0 vdd vdd lock m1_19675_2344# pfet$59
Xpfet$50_4 vdd m1_17703_6956# m1_18496_5840# m1_15755_6960# pfet$50
Xnfet$58_10 m1_12790_7868# vss m1_15618_7156# vss nfet$58
Xpfet$45_7 vdd vdd m1_2446_1478# m1_208_n340# pfet$45
Xnfet$51_6 m1_n940_4493# vss m1_n1212_4493# m1_n1212_4493# m1_n1212_4493# m1_n940_4493#
+ m1_n940_4493# vss m1_n1212_4493# vss nfet$51
Xpfet$50_5 vdd m1_15979_5220# m1_16243_5840# m1_15618_7156# pfet$50
Xnfet$58_11 m1_15979_5220# vss m1_16599_5522# vss nfet$58
Xnfet$58_0 m1_15979_2344# vss m1_16599_2028# vss nfet$58
Xnfet$51_7 m1_3254_4493# vss m1_2982_4493# m1_2982_4493# m1_2982_4493# m1_3254_4493#
+ m1_3254_4493# vss m1_2982_4493# vss nfet$51
Xpfet$50_6 vdd m1_16599_5522# m1_17703_6956# m1_15618_7156# pfet$50
Xpfet$49_10 vdd vdd m1_15618_7156# m1_12790_7868# pfet$49
Xnfet$58_12 m1_15618_7156# vss m1_15755_6960# vss nfet$58
Xnfet$58_1 m1_15618_394# vss m1_15755_n208# vss nfet$58
Xpfet$57_0 vdd vdd m1_n2336_5099# m1_n4030_5270# pfet$57
Xpfet$49_11 vdd vdd m1_16599_5522# m1_15979_5220# pfet$49
Xpfet$50_7 vdd m1_16242_6960# m1_15979_5220# m1_15755_6960# pfet$50
Xnfet$58_13 ref vss m1_16242_6960# vss nfet$58
Xnfet$58_2 m1_n2336_5099# vss m1_16242_n208# vss nfet$58
Xpfet$49_12 vdd vdd m1_16242_6960# ref pfet$49
Xnfet$63_0 m1_19675_2344# vss lock vss nfet$63
Xnfet$56_0 m1_15755_n208# m1_16599_2028# m1_17703_788# vss nfet$56
Xnfet$58_3 m1_17926_34# vss m1_18496_1828# vss nfet$58
Xpfet$49_13 vdd vdd m1_15755_6960# m1_15618_7156# pfet$49
Xnfet$58_4 m1_12790_n340# vss m1_15618_394# vss nfet$58
Xnfet$56_1 m1_15618_394# m1_16242_n208# m1_15979_2344# vss nfet$56
Xnfet$49_0 m1_8596_n340# m1_8596_n340# vss m1_7448_n340# m1_7448_n340# m1_8596_n340#
+ vss m1_7448_n340# m1_7448_n340# m1_7448_n340# m1_8596_n340# m1_7448_n340# m1_7448_n340#
+ m1_8596_n340# vss m1_7448_n340# vss vss nfet$49
Xpfet$55_0 vdd vdd m1_n8022_5099# m1_n10260_7868# pfet$55
Xnfet$58_5 vss vss m1_17215_2028# vss nfet$58
Xnfet$49_1 m1_4402_n340# m1_4402_n340# vss m1_3254_n340# m1_3254_n340# m1_4402_n340#
+ vss m1_3254_n340# m1_3254_n340# m1_3254_n340# m1_4402_n340# m1_3254_n340# m1_3254_n340#
+ m1_4402_n340# vss m1_3254_n340# vss vss nfet$49
Xnfet$56_2 m1_15618_394# m1_17703_788# m1_18496_1828# vss nfet$56
Xpfet$48_0 m1_7448_n340# vdd vdd m1_7448_n340# m1_7176_n340# m1_7176_n340# m1_7448_n340#
+ vdd m1_7176_n340# m1_7176_n340# pfet$48
Xnfet$61_0 m1_n4030_5270# vss m1_n2336_5099# vss nfet$61
Xpfet$55_1 vdd vdd m1_n16410_5099# div pfet$55
.ends

.subckt pfet$85 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=9.75p pd=31.3u as=9.75p ps=31.3u w=15u l=0.5u
.ends

.subckt nfet$91 a_n84_0# a_38_n132# a_138_0# VSUBS
X0 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.5u
.ends

.subckt pfet$86 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=9.75p pd=31.3u as=9.75p ps=31.3u w=15u l=0.5u
.ends

.subckt nfet$92 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$90 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.5u
.ends

.subckt cap_mim$3 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
.ends

.subckt pfet$87 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt CSRVCO_20250823$1 vctrl vosc vdd vss
Xpfet$85_1 vdd vdd m1_n14208_3657# m1_n16019_266# pfet$85
Xnfet$91_0 vss vss vss vss nfet$91
Xpfet$85_2 vdd vdd m1_n13722_3340# m1_n16019_266# pfet$85
Xnfet$91_1 vss vss vss vss nfet$91
Xpfet$85_4 vdd vdd m1_n13236_3035# m1_n16019_266# pfet$85
Xpfet$85_3 vdd m1_n16019_266# vdd m1_n16019_266# pfet$85
Xpfet$85_5 vdd vdd m1_n14693_3963# m1_n16019_266# pfet$85
Xpfet$85_6 vdd vdd m1_n12750_2729# m1_n16019_266# pfet$85
Xpfet$85_7 vdd vdd m1_n15180_4275# m1_n16019_266# pfet$85
Xpfet$85_8 vdd m1_n13236_3035# m1_n9838_266# m1_n10324_266# pfet$85
Xpfet$85_9 vdd m1_n12750_2729# m1_n9352_266# m1_n9838_266# pfet$85
Xpfet$85_10 vdd m1_n14208_3657# m1_n10810_266# m1_n11296_266# pfet$85
Xpfet$85_11 vdd m1_n12264_2422# m1_n11916_1270# m1_n9352_266# pfet$85
Xpfet$85_12 vdd m1_n14693_3963# m1_n11296_266# m1_n11782_266# pfet$85
Xpfet$85_13 vdd m1_n13722_3340# m1_n10324_266# m1_n10810_266# pfet$85
Xpfet$85_14 vdd m1_n15180_4275# m1_n11782_266# m1_n11916_1270# pfet$85
Xpfet$86_0 vdd vdd vdd vdd pfet$86
Xpfet$86_1 vdd vdd vdd vdd pfet$86
Xnfet$92_0 m1_n8380_274# vss vosc vss nfet$92
Xnfet$92_1 m1_n11916_1270# vss m1_n8380_274# vss nfet$92
Xnfet$90_0 m1_n9838_266# m1_n12754_674# m1_n9352_266# vss nfet$90
Xnfet$90_1 vctrl vss m1_n12268_985# vss nfet$90
Xnfet$90_2 vctrl vss m1_n14283_186# vss nfet$90
Xnfet$90_3 vctrl vss m1_n13794_186# vss nfet$90
Xcap_mim$3_0 vss m1_n11296_266# cap_mim$3
Xnfet$90_4 vctrl vss m1_n13240_368# vss nfet$90
Xcap_mim$3_2 vss m1_n10324_266# cap_mim$3
Xcap_mim$3_1 vss m1_n10810_266# cap_mim$3
Xnfet$90_5 vctrl vss m1_n12754_674# vss nfet$90
Xcap_mim$3_3 vss m1_n11916_1270# cap_mim$3
Xnfet$90_6 vctrl m1_n16019_266# vss vss nfet$90
Xnfet$90_7 vctrl vss m1_n15245_186# vss nfet$90
Xcap_mim$3_4 vss m1_n9352_266# cap_mim$3
Xnfet$90_8 vctrl vss m1_n14765_186# vss nfet$90
Xnfet$90_9 m1_n10324_266# m1_n13240_368# m1_n9838_266# vss nfet$90
Xcap_mim$3_5 vss m1_n9838_266# cap_mim$3
Xcap_mim$3_6 vss m1_n11782_266# cap_mim$3
Xnfet$90_10 m1_n9352_266# m1_n12268_985# m1_n11916_1270# vss nfet$90
Xpfet$87_0 vdd vdd vosc m1_n8380_274# pfet$87
Xnfet$90_11 m1_n11916_1270# m1_n15245_186# m1_n11782_266# vss nfet$90
Xpfet$87_1 vdd vdd m1_n8380_274# m1_n11916_1270# pfet$87
Xnfet$90_12 m1_n11782_266# m1_n14765_186# m1_n11296_266# vss nfet$90
Xnfet$90_13 m1_n11296_266# m1_n14283_186# m1_n10810_266# vss nfet$90
Xnfet$90_14 m1_n10810_266# m1_n13794_186# m1_n10324_266# vss nfet$90
Xpfet$85_0 vdd vdd m1_n12264_2422# m1_n16019_266# pfet$85
.ends

.subckt top_level_20250912_nosc i_cp_100u div_def div_prc_s8 div_prc_s7 div_prc_s6
+ div_prc_s5 div_prc_s4 div_prc_s3 div_prc_s2 div_prc_s1 div_prc_s0 div_out div_swc_s0
+ div_swc_s1 div_swc_s2 div_swc_s3 div_swc_s4 div_swc_s5 div_swc_s6 div_swc_s7 div_swc_s8
+ ref ext_pfd_div ext_pfd_ref ext_pfd_up ext_pfd_down mx_pfd_s1 mx_pfd_s0 down cp_s1
+ cp_s2 cp_s3 cp_s4 filter_in filter_out mx_vco_s0 mx_vco_s1 div_rpc_s0 div_rsc_s0
+ div_rsc_s1 div_rpc_s1 div_rsc_s2 div_rpc_s2 div_rsc_s3 div_rsc_s4 div_rsc_s5 div_rsc_s6
+ div_rsc_s7 div_rsc_s8 div_rpc_s3 div_rpc_s4 div_rpc_s5 div_rpc_s6 div_rpc_s7 div_rpc_s8
+ mx_ref_s1 mx_ref_s0 xp_3_1_MUX$5_0/B_1 BIAS$1_0/200n vss vdd xp_3_1_MUX$5_1/B_1
+ div_in ext_vco_out BIAS$1_0/200p2 BIAS$1_0/200p1 up lock out ext_vco_in
Xxp_3_1_MUX$5_2 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX$5_2/OUT_1 xp_3_1_MUX$5_2/C_1
+ xp_3_1_MUX$5_2/B_1 ext_pfd_up xp_3_1_MUX$5
Xxp_3_1_MUX$5_1 mx_vco_s0 mx_vco_s1 vdd vss filter_out xp_3_1_MUX$5_1/C_1 xp_3_1_MUX$5_1/B_1
+ ext_vco_in xp_3_1_MUX$5
Xxp_3_1_MUX$5_3 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX$5_3/OUT_1 xp_3_1_MUX$5_3/C_1
+ xp_3_1_MUX$5_3/B_1 ext_pfd_ref xp_3_1_MUX$5
Xxp_3_1_MUX$5_4 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX$5_4/OUT_1 xp_3_1_MUX$5_4/C_1
+ xp_3_1_MUX$5_4/B_1 ext_pfd_div xp_3_1_MUX$5
Xasc_dual_psd_def_20250809$5_0 vdd vss div_prc_s0 div_prc_s1 div_prc_s2 div_prc_s3
+ div_prc_s4 div_prc_s5 div_prc_s6 div_prc_s7 div_prc_s8 xp_3_1_MUX$5_4/OUT_1 div_swc_s0
+ div_swc_s1 div_swc_s2 div_swc_s3 div_swc_s4 div_swc_s5 div_swc_s6 div_swc_s7 div_swc_s8
+ asc_drive_buffer$5_0/in div_def asc_dual_psd_def_20250809$5
Xxp_3_1_MUX$5_5 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX$5_5/OUT_1 xp_3_1_MUX$5_5/C_1
+ xp_3_1_MUX$5_5/B_1 ext_pfd_down xp_3_1_MUX$5
Xasc_hysteresis_buffer$11_0 vss ref vdd xp_3_1_MUX$6_0/OUT_1 asc_hysteresis_buffer$11
Xasc_drive_buffer$5_0 vss asc_drive_buffer$5_0/in vdd div_in asc_drive_buffer$5
Xasc_drive_buffer$5_1 vss xp_3_1_MUX$5_0/OUT_1 vdd out asc_drive_buffer$5
Xasc_drive_buffer$5_2 vss xp_3_1_MUX$5_4/OUT_1 vdd div_out asc_drive_buffer$5
Xasc_drive_buffer$5_3 vss asc_drive_buffer$5_3/in vdd lock asc_drive_buffer$5
Xasc_drive_buffer$5_4 vss xp_3_1_MUX$5_2/OUT_1 vdd up asc_drive_buffer$5
Xasc_drive_buffer$5_6 vss xp_3_1_MUX$5_5/OUT_1 vdd asc_drive_buffer$5_6/out asc_drive_buffer$5
Xasc_drive_buffer$5_5 vss xp_3_1_MUX$5_5/OUT_1 vdd down asc_drive_buffer$5
Xxp_3_1_MUX$6_0 mx_ref_s0 mx_ref_s1 vdd vss xp_3_1_MUX$6_0/OUT_1 xp_3_1_MUX$6_1/C_1
+ xp_3_1_MUX$6_0/B_1 xp_3_1_MUX$6_0/A_1 xp_3_1_MUX$6
Xxp_3_1_MUX$6_1 mx_ref_s0 mx_ref_s1 vdd vss xp_3_1_MUX$6_1/OUT_1 xp_3_1_MUX$6_1/C_1
+ xp_3_1_MUX$6_1/B_1 xp_3_1_MUX$6_1/A_1 xp_3_1_MUX$6
Xasc_dual_psd_def_20250809$6_0 vdd vss div_rpc_s0 div_rpc_s1 div_rpc_s2 div_rpc_s3
+ div_rpc_s4 div_rpc_s5 div_rpc_s6 div_rpc_s7 div_rpc_s8 xp_3_1_MUX$6_1/B_1 div_rsc_s0
+ div_rsc_s1 div_rsc_s2 div_rsc_s3 div_rsc_s4 div_rsc_s5 div_rsc_s6 div_rsc_s7 div_rsc_s8
+ xp_3_1_MUX$6_0/B_1 vss asc_dual_psd_def_20250809$6
Xasc_drive_buffer$6_0 vss xp_3_1_MUX$5_0/OUT_1 vdd asc_drive_buffer$5_0/in asc_drive_buffer$6
Xasc_hysteresis_buffer$10_0 vss xp_3_1_MUX$6_1/OUT_1 vdd xp_3_1_MUX$5_3/OUT_1 asc_hysteresis_buffer$10
Xxp_programmable_basic_pump$1_0 asc_drive_buffer_up$1_0/out vdd cp_s1 cp_s2 cp_s3
+ cp_s4 asc_drive_buffer$5_6/out filter_in BIAS$1_0/100n vss xp_programmable_basic_pump$1
Xasc_PFD_DFF_20250831$1_0 vss xp_3_1_MUX$5_3/C_1 xp_3_1_MUX$5_5/C_1 xp_3_1_MUX$5_2/C_1
+ vdd xp_3_1_MUX$5_4/C_1 asc_PFD_DFF_20250831$1
Xasc_PFD_DFF_20250831$1_1 vss xp_3_1_MUX$5_3/B_1 xp_3_1_MUX$5_2/B_1 xp_3_1_MUX$5_5/B_1
+ vdd xp_3_1_MUX$5_4/B_1 asc_PFD_DFF_20250831$1
Xasc_drive_buffer_up$1_0 vss asc_drive_buffer_up$1_0/out xp_3_1_MUX$5_2/OUT_1 vdd
+ asc_drive_buffer_up$1
XBIAS$1_0 vdd vss BIAS$1_0/100n BIAS$1_0/200n i_cp_100u BIAS$1_0/200p1 BIAS$1_0/200p2
+ BIAS$1
Xasc_lock_detector_20250826$1_0 xp_3_1_MUX$5_3/OUT_1 vdd xp_3_1_MUX$5_4/OUT_1 vss
+ asc_drive_buffer$5_3/in asc_lock_detector_20250826$1
XCSRVCO_20250823$1_0 xp_3_1_MUX$5_1/C_1 xp_3_1_MUX$5_0/C_1 vdd vss CSRVCO_20250823$1
Xxp_3_1_MUX$5_0 mx_vco_s0 mx_vco_s1 vdd vss xp_3_1_MUX$5_0/OUT_1 xp_3_1_MUX$5_0/C_1
+ xp_3_1_MUX$5_0/B_1 ext_vco_out xp_3_1_MUX$5
.ends

.subckt pfet$102 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=0.8125p pd=3.8u as=0.325p ps=1.77u w=1.25u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.325p pd=1.77u as=0.8125p ps=3.8u w=1.25u l=0.5u
.ends

.subckt pfet$101 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# w_n180_n88# a_1262_n60# a_38_n60# a_n92_0# a_1058_n60# a_854_n60# a_342_0#
+ a_138_0# a_650_n60# a_1362_0#
X0 a_1362_0# a_1262_n60# a_1158_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X1 a_954_0# a_854_n60# a_750_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X2 a_1566_0# a_1466_n60# a_1362_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.5u
X3 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X4 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X5 a_1158_0# a_1058_n60# a_954_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X6 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.5u
X7 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
.ends

.subckt nfet$110 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$107 a_750_0# a_546_0# a_446_n132# a_n84_0# a_650_n132# a_38_n132# a_342_0#
+ a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.5u
X1 a_546_0# a_446_n132# a_342_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.5u
X2 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.5u
X3 a_750_0# a_650_n132# a_546_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.5u
.ends

.subckt nfet$111 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.5u
.ends

.subckt nfet$106 a_30_n132# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt cap_mim$4 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=50u c_length=100u
.ends

.subckt nfet$108 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$105 a_750_0# a_546_0# a_446_n60# a_242_n60# w_n180_n88# a_38_n60# a_n92_0#
+ a_342_0# a_138_0# a_650_n60#
X0 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X2 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.5u
.ends

.subckt pfet$100 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
.ends

.subckt pfet$99 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_348_n136# a_414_0# a_n92_0#
+ a_94_0# a_574_0# a_508_n136#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_n136# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_n136# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$104 a_254_0# a_30_n132# a_n84_0# a_94_0# a_190_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt nfet$105 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt OTAforChargePump$1 vdd vss out iref inn inp
Xpfet$100_0 m1_n400_n914# m1_n400_n914# m1_n400_n914# vdd m1_n400_n914# m1_n400_n914#
+ pfet$100
Xpfet$100_1 m1_n400_n914# m1_n400_n914# m1_n400_n914# vdd m1_n400_n914# m1_n400_n914#
+ pfet$100
Xpfet$100_2 vdd vdd vdd vdd vdd vdd pfet$100
Xpfet$100_3 vdd vdd vdd vdd vdd vdd pfet$100
Xpfet$100_5 vdd vdd vdd vdd vdd vdd pfet$100
Xpfet$100_4 vdd vdd vdd vdd vdd vdd pfet$100
Xpfet$99_0 inn m1_n400_n914# inn vdd inn out m1_n400_n914# out m1_n400_n914# inn pfet$99
Xpfet$99_1 inp m1_n400_n914# inp vdd inp m1_116_n1334# m1_n400_n914# m1_116_n1334#
+ m1_n400_n914# inp pfet$99
Xpfet$99_2 iref vdd iref vdd iref iref vdd iref vdd iref pfet$99
Xpfet$99_3 iref vdd iref vdd iref m1_n400_n914# vdd m1_n400_n914# vdd iref pfet$99
Xpfet$99_4 iref vdd iref vdd iref m1_n400_n914# vdd m1_n400_n914# vdd iref pfet$99
Xpfet$99_6 iref vdd iref vdd iref iref vdd iref vdd iref pfet$99
Xpfet$99_5 iref vdd iref vdd iref iref vdd iref vdd iref pfet$99
Xpfet$99_11 iref vdd iref vdd iref m1_n400_n914# vdd m1_n400_n914# vdd iref pfet$99
Xpfet$99_10 iref vdd iref vdd iref iref vdd iref vdd iref pfet$99
Xpfet$99_7 iref vdd iref vdd iref m1_n400_n914# vdd m1_n400_n914# vdd iref pfet$99
Xpfet$99_8 inp m1_n400_n914# inp vdd inp m1_116_n1334# m1_n400_n914# m1_116_n1334#
+ m1_n400_n914# inp pfet$99
Xpfet$99_9 inn m1_n400_n914# inn vdd inn out m1_n400_n914# out m1_n400_n914# inn pfet$99
Xnfet$104_1 vss m1_116_n1334# vss m1_116_n1334# m1_116_n1334# vss nfet$104
Xnfet$104_0 vss m1_116_n1334# vss out m1_116_n1334# vss nfet$104
Xnfet$104_2 vss m1_116_n1334# vss m1_116_n1334# m1_116_n1334# vss nfet$104
Xnfet$104_3 vss m1_116_n1334# vss out m1_116_n1334# vss nfet$104
Xnfet$105_0 vss vss vss vss vss vss vss vss vss vss nfet$105
Xnfet$105_1 vss vss vss vss vss vss vss vss vss vss nfet$105
.ends

.subckt pfet$103 a_28_460# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_460# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt nfet$109 a_750_0# a_546_0# a_446_n132# a_n84_0# a_650_n132# a_38_n132# a_342_0#
+ a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_546_0# a_446_n132# a_342_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X2 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
X3 a_750_0# a_650_n132# a_546_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt pfet$106 a_1054_0# a_734_0# a_828_n136# a_28_n136# a_254_0# a_894_0# a_188_n136#
+ a_988_n136# w_n180_n88# a_348_n136# a_1214_0# a_1148_n136# a_414_0# a_n92_0# a_94_0#
+ a_574_0# a_508_n136# a_668_n136#
X0 a_1214_0# a_1148_n136# a_1054_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_734_0# a_668_n136# a_574_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X3 a_574_0# a_508_n136# a_414_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X4 a_1054_0# a_988_n136# a_894_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X5 a_894_0# a_828_n136# a_734_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X6 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X7 a_414_0# a_348_n136# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt ppolyf_u_resistor$1 a_4000_0# a_n376_0# a_n132_0#
X0 a_n132_0# a_4000_0# a_n376_0# ppolyf_u r_width=1u r_length=20u
.ends

.subckt pfet$104 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$112 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt PCP1248X$1 vdd s3 s2 s1 s0 vin iref200u out up down vss
Xpfet$102_3 vdd vdd vdd m1_n1751_n2187# m1_n1751_n2187# m1_n1751_n2187# pfet$102
Xpfet$101_14 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$101
Xpfet$101_25 vdd vdd m1_1671_n1319# m1_1137_12199# m1_1137_12199# vdd m1_1671_n1319#
+ m1_1137_12199# vdd m1_1137_12199# m1_1137_12199# vdd m1_1137_12199# m1_1137_12199#
+ vdd m1_1671_n1319# m1_1137_12199# m1_1671_n1319# pfet$101
Xnfet$110_2 s1 vss m1_n1311_12403# vss nfet$110
Xnfet$107_8 m1_13543_n1758# m1_15911_n1318# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15911_n1318# m1_9963_14448# vss nfet$107
Xpfet$102_4 vdd vdd vdd m1_9963_14448# m1_n1751_n2187# m1_n1751_n2187# pfet$102
Xnfet$110_3 s0 vss m1_n539_12403# vss nfet$110
Xpfet$101_15 m1_n2925_n36# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187#
+ m1_1671_n1319# pfet$101
Xpfet$101_26 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$101
Xnfet$107_9 m1_13543_n1758# m1_15911_n1318# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15911_n1318# m1_9963_14448# vss nfet$107
Xpfet$102_5 vdd vdd vdd vdd vdd vdd pfet$102
Xpfet$101_16 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ pfet$101
Xpfet$101_27 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$101
Xnfet$111_10 vss vss vss vss vss vss nfet$111
Xnfet$106_10 m1_n2855_12403# m1_14137_3830# vss vss nfet$106
Xpfet$101_17 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$101
Xpfet$101_28 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$101
Xnfet$106_11 s3 OTAforChargePump$1_0/out m1_14137_3830# vss nfet$106
Xnfet$111_11 vss vss vss vss vss vss nfet$111
Xcap_mim$4_0 m1_n1751_n2187# vdd cap_mim$4
Xpfet$101_18 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$101
Xpfet$101_29 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ pfet$101
Xcap_mim$4_1 vss m1_9963_14448# cap_mim$4
Xpfet$101_19 m1_n2925_n36# m1_n2925_n36# m1_n25_493# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n25_493# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36#
+ m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n25_493# m1_n1751_n2187# m1_n25_493#
+ pfet$101
Xcap_mim$4_2 vss OTAforChargePump$1_0/out cap_mim$4
Xnfet$108_0 vss vss vss vss vss vss nfet$108
Xpfet$105_10 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$105
Xnfet$108_1 vss vss vss vss vss vss nfet$108
Xpfet$105_11 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$105
Xpfet$105_0 m1_n47_11059# m1_n47_11059# m1_n47_11059# m1_n47_11059# vdd m1_n47_11059#
+ m1_n47_11059# m1_n47_11059# m1_n47_11059# m1_n47_11059# pfet$105
Xnfet$108_2 vss m1_9963_14448# vss m1_9963_14448# m1_9963_14448# vss nfet$108
Xpfet$105_1 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$105
XOTAforChargePump$1_0 vdd vss OTAforChargePump$1_0/out iref200u vin OTAforChargePump$1_0/inp
+ OTAforChargePump$1
Xnfet$106_0 s0 m1_n47_11059# m1_1641_5849# vss nfet$106
Xpfet$105_2 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$105
Xnfet$107_30 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$107
Xpfet$105_3 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$105
Xnfet$106_1 s1 m1_n47_11059# m1_n91_6229# vss nfet$106
Xpfet$103_0 s0 vdd m1_1641_5849# vdd pfet$103
Xnfet$107_20 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$107
Xnfet$106_2 s3 m1_n47_11059# m1_n1771_4009# vss nfet$106
Xnfet$107_31 m1_n47_11059# m1_14015_1164# m1_9963_14448# m1_n47_11059# m1_9963_14448#
+ m1_9963_14448# m1_n47_11059# m1_14015_1164# m1_9963_14448# vss nfet$107
Xpfet$105_4 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$105
Xpfet$103_1 s3 vdd m1_n1771_4009# vdd pfet$103
Xnfet$111_0 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$111
Xnfet$107_21 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$107
Xnfet$107_32 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$107
Xnfet$107_10 m1_13543_n1758# m1_15911_n1318# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15911_n1318# m1_9963_14448# vss nfet$107
Xnfet$106_3 s2 m1_n47_11059# m1_1137_12199# vss nfet$106
Xpfet$105_5 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$105
Xpfet$103_2 m1_n1311_12403# vdd m1_n47_11059# m1_n91_6229# pfet$103
Xnfet$111_1 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$111
Xnfet$106_4 m1_n539_12403# m1_16753_5552# vss vss nfet$106
Xnfet$107_22 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$107
Xnfet$107_33 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$107
Xnfet$107_11 m1_13543_n1758# m1_15039_784# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15039_784# m1_9963_14448# vss nfet$107
Xpfet$105_6 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$105
Xpfet$103_3 m1_n2083_12403# vdd m1_n47_11059# m1_1137_12199# pfet$103
Xnfet$111_2 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$111
Xpfet$101_0 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$101
Xnfet$107_34 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$107
Xnfet$107_23 vss m1_15039_784# m1_15009_5932# vss m1_15009_5932# m1_15009_5932# vss
+ m1_15039_784# m1_15009_5932# vss nfet$107
Xnfet$107_12 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$107
Xnfet$106_5 s0 OTAforChargePump$1_0/out m1_16753_5552# vss nfet$106
Xpfet$105_7 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$105
Xpfet$103_4 m1_n2855_12403# vdd m1_n47_11059# m1_n1771_4009# pfet$103
Xnfet$111_3 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$111
Xpfet$101_1 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$101
Xnfet$107_24 vss vss vss vss vss vss vss vss vss vss nfet$107
Xnfet$107_35 vss m1_14015_1164# OTAforChargePump$1_0/out vss OTAforChargePump$1_0/out
+ OTAforChargePump$1_0/out vss m1_14015_1164# OTAforChargePump$1_0/out vss nfet$107
Xnfet$107_13 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$107
Xnfet$106_6 m1_n1311_12403# m1_15009_5932# vss vss nfet$106
Xpfet$105_8 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$105
Xpfet$103_5 s1 vdd m1_n91_6229# vdd pfet$103
Xnfet$111_4 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$111
Xpfet$101_2 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$101
Xnfet$107_36 OTAforChargePump$1_0/inp m1_9475_12045# m1_9963_14448# OTAforChargePump$1_0/inp
+ m1_9963_14448# m1_9963_14448# OTAforChargePump$1_0/inp m1_9475_12045# m1_9963_14448#
+ vss nfet$107
Xnfet$107_25 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$107
Xnfet$107_14 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$107
Xnfet$106_7 s1 OTAforChargePump$1_0/out m1_15009_5932# vss nfet$106
Xpfet$105_9 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$105
Xpfet$103_6 s2 vdd m1_1137_12199# vdd pfet$103
Xnfet$111_5 m1_n47_11059# m1_n47_11059# m1_n47_11059# m1_n47_11059# m1_n47_11059#
+ vss nfet$111
Xpfet$101_3 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$101
Xnfet$107_26 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$107
Xnfet$107_15 vss vss vss vss vss vss vss vss vss vss nfet$107
Xnfet$106_8 m1_n2083_12403# m1_15881_3450# vss vss nfet$106
Xnfet$111_6 vss vss vss vss vss vss nfet$111
Xpfet$103_7 m1_n539_12403# vdd m1_n47_11059# m1_1641_5849# pfet$103
Xpfet$103_10 m1_n2083_12403# vdd OTAforChargePump$1_0/out m1_15881_3450# pfet$103
Xpfet$101_4 m1_n2925_n36# m1_n2925_n36# m1_n25_493# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n25_493# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36#
+ m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n25_493# m1_n1751_n2187# m1_n25_493#
+ pfet$101
Xnfet$106_9 s2 OTAforChargePump$1_0/out m1_15881_3450# vss nfet$106
Xnfet$107_27 vss m1_15911_n1318# m1_15881_3450# vss m1_15881_3450# m1_15881_3450#
+ vss m1_15911_n1318# m1_15881_3450# vss nfet$107
Xnfet$107_16 vss m1_16783_404# m1_16753_5552# vss m1_16753_5552# m1_16753_5552# vss
+ m1_16783_404# m1_16753_5552# vss nfet$107
Xpfet$103_8 m1_n539_12403# vdd OTAforChargePump$1_0/out m1_16753_5552# pfet$103
Xnfet$111_7 vss vss vss vss vss vss nfet$111
Xpfet$103_11 m1_n2855_12403# vdd OTAforChargePump$1_0/out m1_14137_3830# pfet$103
Xpfet$101_5 m1_n47_11059# m1_n47_11059# m1_6759_7857# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n47_11059# m1_6759_7857# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n47_11059# m1_n1751_n2187# m1_n1751_n2187# m1_n47_11059# m1_6759_7857# m1_n1751_n2187#
+ m1_6759_7857# pfet$101
Xnfet$107_28 vss m1_15911_n1318# m1_15881_3450# vss m1_15881_3450# m1_15881_3450#
+ vss m1_15911_n1318# m1_15881_3450# vss nfet$107
Xnfet$107_17 vss m1_15039_784# m1_15009_5932# vss m1_15009_5932# m1_15009_5932# vss
+ m1_15039_784# m1_15009_5932# vss nfet$107
Xnfet$111_8 vss vss vss vss vss vss nfet$111
Xpfet$103_9 m1_n1311_12403# vdd OTAforChargePump$1_0/out m1_15009_5932# pfet$103
Xpfet$101_6 vdd vdd m1_6759_7857# m1_n47_11059# m1_n47_11059# vdd m1_6759_7857# m1_n47_11059#
+ vdd m1_n47_11059# m1_n47_11059# vdd m1_n47_11059# m1_n47_11059# vdd m1_6759_7857#
+ m1_n47_11059# m1_6759_7857# pfet$101
Xnfet$107_29 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$107
Xnfet$107_18 vss m1_15911_n1318# m1_15881_3450# vss m1_15881_3450# m1_15881_3450#
+ vss m1_15911_n1318# m1_15881_3450# vss nfet$107
Xnfet$111_9 vss vss vss vss vss vss nfet$111
Xpfet$101_7 vdd vdd m1_n25_493# m1_n91_6229# m1_n91_6229# vdd m1_n25_493# m1_n91_6229#
+ vdd m1_n91_6229# m1_n91_6229# vdd m1_n91_6229# m1_n91_6229# vdd m1_n25_493# m1_n91_6229#
+ m1_n25_493# pfet$101
Xnfet$107_19 vss m1_15911_n1318# m1_15881_3450# vss m1_15881_3450# m1_15881_3450#
+ vss m1_15911_n1318# m1_15881_3450# vss nfet$107
Xpfet$101_8 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$101
Xnfet$109_0 vss m1_9475_12045# OTAforChargePump$1_0/out vss OTAforChargePump$1_0/out
+ OTAforChargePump$1_0/out vss m1_9475_12045# OTAforChargePump$1_0/out vss nfet$109
Xpfet$101_9 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$101
Xnfet$109_1 vss m1_n1751_n2187# OTAforChargePump$1_0/out vss OTAforChargePump$1_0/out
+ OTAforChargePump$1_0/out vss m1_n1751_n2187# OTAforChargePump$1_0/out vss nfet$109
Xpfet$106_0 m1_n2925_n36# m1_n2925_n36# up up out out up up vdd up out up m1_n2925_n36#
+ out m1_n2925_n36# out up up pfet$106
Xnfet$109_2 vss m1_9475_12045# OTAforChargePump$1_0/out vss OTAforChargePump$1_0/out
+ OTAforChargePump$1_0/out vss m1_9475_12045# OTAforChargePump$1_0/out vss nfet$109
Xnfet$109_3 vss m1_n1751_n2187# OTAforChargePump$1_0/out vss OTAforChargePump$1_0/out
+ OTAforChargePump$1_0/out vss m1_n1751_n2187# OTAforChargePump$1_0/out vss nfet$109
Xppolyf_u_resistor$1_0 m1_3630_13790# vss m1_n502_13390# ppolyf_u_resistor$1
Xnfet$107_0 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$107
Xnfet$107_1 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$107
Xpfet$104_0 vdd vdd m1_n2855_12403# s3 pfet$104
Xppolyf_u_resistor$1_1 OTAforChargePump$1_0/inp vss m1_n502_13390# ppolyf_u_resistor$1
Xpfet$101_30 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ pfet$101
Xppolyf_u_resistor$1_2 m1_3630_14590# vss m1_n502_14190# ppolyf_u_resistor$1
Xnfet$112_0 down out m1_13543_n1758# down out m1_13543_n1758# down out down vss nfet$112
Xnfet$107_2 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$107
Xpfet$104_1 vdd vdd m1_n2083_12403# s2 pfet$104
Xpfet$101_31 m1_n2925_n36# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187#
+ m1_1671_n1319# pfet$101
Xpfet$101_20 m1_n2925_n36# m1_n2925_n36# m1_1671_873# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_873# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36#
+ m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_873# m1_n1751_n2187# m1_1671_873#
+ pfet$101
Xnfet$107_3 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# vss nfet$107
Xpfet$104_2 vdd vdd m1_n539_12403# s0 pfet$104
Xppolyf_u_resistor$1_3 m1_3630_13790# vss m1_n502_14190# ppolyf_u_resistor$1
Xpfet$101_10 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$101
Xpfet$101_32 m1_n2925_n36# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187#
+ m1_1671_n1319# pfet$101
Xpfet$101_21 vdd vdd m1_1671_873# m1_1641_5849# m1_1641_5849# vdd m1_1671_873# m1_1641_5849#
+ vdd m1_1641_5849# m1_1641_5849# vdd m1_1641_5849# m1_1641_5849# vdd m1_1671_873#
+ m1_1641_5849# m1_1671_873# pfet$101
Xppolyf_u_resistor$1_4 m1_3630_14590# vss m1_n502_14990# ppolyf_u_resistor$1
Xnfet$107_4 m1_13543_n1758# m1_15039_784# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15039_784# m1_9963_14448# vss nfet$107
Xpfet$102_0 vdd vdd vdd vdd vdd vdd pfet$102
Xpfet$104_3 vdd vdd m1_n1311_12403# s1 pfet$104
Xpfet$101_11 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$101
Xpfet$101_22 vdd vdd m1_1671_n1319# m1_1137_12199# m1_1137_12199# vdd m1_1671_n1319#
+ m1_1137_12199# vdd m1_1137_12199# m1_1137_12199# vdd m1_1137_12199# m1_1137_12199#
+ vdd m1_1671_n1319# m1_1137_12199# m1_1671_n1319# pfet$101
Xpfet$101_33 vdd vdd m1_1671_n1319# m1_1137_12199# m1_1137_12199# vdd m1_1671_n1319#
+ m1_1137_12199# vdd m1_1137_12199# m1_1137_12199# vdd m1_1137_12199# m1_1137_12199#
+ vdd m1_1671_n1319# m1_1137_12199# m1_1671_n1319# pfet$101
Xnfet$107_5 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# vss nfet$107
Xppolyf_u_resistor$1_5 vdd vss m1_n502_14990# ppolyf_u_resistor$1
Xpfet$102_1 vdd vdd vdd m1_n1751_n2187# m1_n1751_n2187# m1_n1751_n2187# pfet$102
Xpfet$101_12 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$101
Xpfet$101_23 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$101
Xpfet$101_34 vdd vdd m1_1671_n1319# m1_1137_12199# m1_1137_12199# vdd m1_1671_n1319#
+ m1_1137_12199# vdd m1_1137_12199# m1_1137_12199# vdd m1_1137_12199# m1_1137_12199#
+ vdd m1_1671_n1319# m1_1137_12199# m1_1671_n1319# pfet$101
Xnfet$110_0 s3 vss m1_n2855_12403# vss nfet$110
Xnfet$107_6 m1_13543_n1758# m1_16783_404# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_16783_404# m1_9963_14448# vss nfet$107
Xpfet$102_2 vdd vdd vdd m1_9963_14448# m1_n1751_n2187# m1_n1751_n2187# pfet$102
Xnfet$110_1 s2 vss m1_n2083_12403# vss nfet$110
Xpfet$101_13 m1_n2925_n36# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187#
+ m1_1671_n1319# pfet$101
Xpfet$101_24 vdd vdd m1_n25_493# m1_n91_6229# m1_n91_6229# vdd m1_n25_493# m1_n91_6229#
+ vdd m1_n91_6229# m1_n91_6229# vdd m1_n91_6229# m1_n91_6229# vdd m1_n25_493# m1_n91_6229#
+ m1_n25_493# pfet$101
Xpfet$101_35 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ pfet$101
Xnfet$107_7 m1_13543_n1758# m1_15911_n1318# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15911_n1318# m1_9963_14448# vss nfet$107
.ends

.subckt pfet$116 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt pfet$107 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt nfet$113 a_n84_0# a_94_0# a_30_160# VSUBS
X0 a_94_0# a_30_160# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.28u
.ends

.subckt SRLATCH vdd vss q qb s r
Xpfet$107_0 r vdd m1_818_875# qb pfet$107
Xpfet$107_1 q vdd vdd m1_818_875# pfet$107
Xpfet$107_2 s vdd m1_50_875# vdd pfet$107
Xpfet$107_3 qb vdd q m1_50_875# pfet$107
Xnfet$113_0 vss qb r vss nfet$113
Xnfet$113_1 vss qb q vss nfet$113
Xnfet$113_3 q vss qb vss nfet$113
Xnfet$113_2 q vss s vss nfet$113
.ends

.subckt ppolyf_u_resistor$2 a_n376_0# a_4200_0# a_n132_0#
X0 a_n132_0# a_4200_0# a_n376_0# ppolyf_u r_width=1u r_length=21u
.ends

.subckt pfet$114 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=2.6p pd=9.3u as=2.6p ps=9.3u w=4u l=0.28u
.ends

.subckt nfet$122 a_30_n132# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$115 a_28_460# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_460# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt nfet$121 a_n84_0# a_94_0# a_30_460# VSUBS
X0 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt SCHMITT$6 VDD VSS IN OUT
Xpfet$114_0 IN VDD m1_596_1544# OUT pfet$114
Xpfet$114_1 IN VDD VDD m1_596_1544# pfet$114
Xnfet$122_0 OUT m1_592_402# VDD VSS nfet$122
Xpfet$115_0 OUT VDD m1_596_1544# VSS pfet$115
Xnfet$121_0 m1_592_402# OUT IN VSS nfet$121
Xnfet$121_1 VSS m1_592_402# IN VSS nfet$121
.ends

.subckt cap_mim$5 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=60u c_length=100u
.ends

.subckt nfet$123 a_30_260# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_260# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$109 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
.ends

.subckt nfet$117 a_n84_0# a_94_0# a_30_460# VSUBS
X0 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt nfet$115 a_1054_0# a_734_0# a_254_0# a_350_460# a_830_460# a_894_0# a_990_460#
+ a_1214_0# a_414_0# a_n84_0# a_94_0# a_510_460# a_190_460# a_574_0# a_670_460# a_1150_460#
+ a_30_460# VSUBS
X0 a_734_0# a_670_460# a_574_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_574_0# a_510_460# a_414_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X3 a_1054_0# a_990_460# a_894_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X4 a_894_0# a_830_460# a_734_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X5 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X6 a_414_0# a_350_460# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X7 a_1214_0# a_1150_460# a_1054_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt pfet$110 a_254_0# a_348_560# w_n180_n88# a_414_0# a_n92_0# a_94_0# a_574_0#
+ a_508_560# a_188_560# a_28_560#
X0 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt pfet$108 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_348_n136# a_414_0#
+ a_n92_0# a_94_0# a_574_0# a_508_n136#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_n136# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_n136# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$116 a_254_0# a_350_460# a_414_0# a_n84_0# a_94_0# a_510_460# a_190_460#
+ a_574_0# a_30_460# VSUBS
X0 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_460# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_460# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt nfet$114 a_254_0# a_n84_0# a_94_0# a_190_460# a_30_460# VSUBS
X0 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt Ncomparator$1 iref vss vdd out inn inp
Xpfet$109_0 vdd vdd vdd vdd vdd vdd pfet$109
Xpfet$109_1 vdd vdd vdd vdd vdd vdd pfet$109
Xnfet$117_0 vss vss vss vss nfet$117
Xpfet$109_2 vdd vdd vdd vdd vdd vdd pfet$109
Xnfet$117_1 vss vss vss vss nfet$117
Xpfet$109_3 vdd vdd vdd vdd vdd vdd pfet$109
Xnfet$115_0 out out vss iref iref vss iref vss out vss out iref iref vss iref iref
+ iref vss nfet$115
Xpfet$110_0 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$110
Xpfet$110_1 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$110
Xpfet$110_2 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$110
Xpfet$110_3 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$110
Xpfet$108_0 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_570_1653# vdd m1_570_1653#
+ vdd m1_1242_549# pfet$108
Xpfet$108_2 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_570_1653# vdd m1_570_1653#
+ vdd m1_1242_549# pfet$108
Xpfet$108_1 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_1242_549# vdd m1_1242_549#
+ vdd m1_1242_549# pfet$108
Xnfet$116_1 vss iref iref vss iref iref iref vss iref vss nfet$116
Xnfet$116_0 vss iref m1_506_n191# vss m1_506_n191# iref iref vss iref vss nfet$116
Xpfet$108_3 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_1242_549# vdd m1_1242_549#
+ vdd m1_1242_549# pfet$108
Xnfet$116_2 m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191#
+ m1_506_n191# m1_506_n191# m1_506_n191# vss nfet$116
Xnfet$116_3 m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191#
+ m1_506_n191# m1_506_n191# m1_506_n191# vss nfet$116
Xnfet$114_0 m1_506_n191# m1_506_n191# m1_570_1653# inp inp vss nfet$114
Xnfet$116_4 vss iref iref vss iref iref iref vss iref vss nfet$116
Xnfet$114_1 m1_506_n191# m1_506_n191# m1_1242_549# inn inn vss nfet$114
Xnfet$114_2 m1_506_n191# m1_506_n191# m1_570_1653# inp inp vss nfet$114
Xnfet$116_5 vss iref m1_506_n191# vss m1_506_n191# iref iref vss iref vss nfet$116
Xnfet$114_3 m1_506_n191# m1_506_n191# m1_1242_549# inn inn vss nfet$114
.ends

.subckt pfet$112 a_254_0# a_348_560# w_n180_n88# a_414_0# a_n92_0# a_94_0# a_574_0#
+ a_508_560# a_188_560# a_28_560#
X0 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$119 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt nfet$120 a_254_0# a_n84_0# a_94_0# a_190_460# a_30_460# VSUBS
X0 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt nfet$118 a_1054_0# a_734_0# a_510_n132# a_254_0# a_894_0# a_670_n132# a_1214_0#
+ a_830_n132# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132# a_574_0# a_990_n132#
+ a_350_n132# a_1150_n132# VSUBS
X0 a_734_0# a_670_n132# a_574_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X3 a_1054_0# a_990_n132# a_894_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X4 a_894_0# a_830_n132# a_734_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X5 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X6 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X7 a_1214_0# a_1150_n132# a_1054_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt pfet$113 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=1.625p ps=6.3u w=2.5u l=0.28u
.ends

.subckt pfet$111 a_1054_0# a_734_0# a_254_0# a_894_0# a_348_560# a_828_560# a_988_560#
+ w_n180_n88# a_1214_0# a_414_0# a_n92_0# a_94_0# a_574_0# a_508_560# a_188_560# a_668_560#
+ a_1148_560# a_28_560#
X0 a_1214_0# a_1148_560# a_1054_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_734_0# a_668_560# a_574_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X3 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X4 a_1054_0# a_988_560# a_894_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X5 a_894_0# a_828_560# a_734_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X6 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X7 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt Pcomparator$1 vss vdd out iref inn inp
Xpfet$112_13 m1_2779_n1752# inp vdd m1_5539_n2811# m1_2779_n1752# m1_5539_n2811# m1_2779_n1752#
+ inp inp inp pfet$112
Xnfet$119_0 vss vss vss vss vss vss vss vss vss vss nfet$119
Xnfet$119_1 vss vss vss vss vss vss vss vss vss vss nfet$119
Xpfet$112_0 m1_2779_n1752# inp vdd m1_5539_n2811# m1_2779_n1752# m1_5539_n2811# m1_2779_n1752#
+ inp inp inp pfet$112
Xpfet$112_1 m1_2779_n1752# m1_2779_n1752# vdd m1_2779_n1752# m1_2779_n1752# m1_2779_n1752#
+ m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# pfet$112
Xnfet$120_0 vss vss m1_3615_n1223# m1_3615_n1223# m1_3615_n1223# vss nfet$120
Xpfet$112_2 m1_2779_n1752# inn vdd m1_3615_n1223# m1_2779_n1752# m1_3615_n1223# m1_2779_n1752#
+ inn inn inn pfet$112
Xnfet$120_1 vss vss m1_5539_n2811# m1_3615_n1223# m1_3615_n1223# vss nfet$120
Xpfet$112_3 m1_2779_n1752# m1_2779_n1752# vdd m1_2779_n1752# m1_2779_n1752# m1_2779_n1752#
+ m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# pfet$112
Xnfet$120_2 vss vss m1_5539_n2811# m1_3615_n1223# m1_3615_n1223# vss nfet$120
Xpfet$112_4 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$112
Xnfet$120_3 vss vss m1_3615_n1223# m1_3615_n1223# m1_3615_n1223# vss nfet$120
Xpfet$112_6 vdd iref vdd iref vdd iref vdd iref iref iref pfet$112
Xpfet$112_5 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$112
Xpfet$112_7 vdd iref vdd iref vdd iref vdd iref iref iref pfet$112
Xpfet$112_8 vdd iref vdd iref vdd iref vdd iref iref iref pfet$112
Xpfet$112_9 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$112
Xnfet$118_0 out out m1_5539_n2811# vss vss m1_5539_n2811# vss m1_5539_n2811# out m1_5539_n2811#
+ vss out m1_5539_n2811# vss m1_5539_n2811# m1_5539_n2811# m1_5539_n2811# vss nfet$118
Xpfet$113_0 vdd vdd vdd vdd pfet$113
Xpfet$113_2 vdd vdd vdd vdd pfet$113
Xpfet$113_1 vdd vdd vdd vdd pfet$113
Xpfet$111_0 out out vdd vdd iref iref iref vdd vdd out vdd out vdd iref iref iref
+ iref iref pfet$111
Xpfet$113_3 vdd vdd vdd vdd pfet$113
Xpfet$111_1 out out vdd vdd iref iref iref vdd vdd out vdd out vdd iref iref iref
+ iref iref pfet$111
Xpfet$112_10 vdd iref vdd iref vdd iref vdd iref iref iref pfet$112
Xpfet$112_11 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$112
Xpfet$112_12 m1_2779_n1752# inn vdd m1_3615_n1223# m1_2779_n1752# m1_3615_n1223# m1_2779_n1752#
+ inn inn inn pfet$112
.ends

.subckt VCOfinal s3 s0 s1 s2 iref200 fout foutb irefn irefp vin vss vdd a_11641_n18839#
XPCP1248X$1_0 vdd s3 s2 s1 s0 vin iref200 PCP1248X$1_0/out PCP1248X$1_0/up SRLATCH_0/qb
+ vss PCP1248X$1
Xpfet$116_0 SRLATCH_0/q vdd vdd PCP1248X$1_0/up pfet$116
Xpfet$116_1 SCHMITT$6_0/OUT vdd vdd foutb pfet$116
Xpfet$116_2 SCHMITT$6_1/OUT vdd vdd fout pfet$116
XSRLATCH_0 vdd vss SRLATCH_0/q SRLATCH_0/qb SRLATCH_0/s SRLATCH_0/r SRLATCH
Xppolyf_u_resistor$2_0 vss vss Pcomparator$1_0/inp ppolyf_u_resistor$2
Xppolyf_u_resistor$2_1 vss m1_13996_n13334# Ncomparator$1_0/inn ppolyf_u_resistor$2
Xppolyf_u_resistor$2_2 vss m1_13996_n13334# Pcomparator$1_0/inp ppolyf_u_resistor$2
XSCHMITT$6_1 vdd vss SRLATCH_0/q SCHMITT$6_1/OUT SCHMITT$6
XSCHMITT$6_0 vdd vss SRLATCH_0/qb SCHMITT$6_0/OUT SCHMITT$6
Xppolyf_u_resistor$2_3 vss vdd Ncomparator$1_0/inn ppolyf_u_resistor$2
Xcap_mim$5_0 vss PCP1248X$1_0/out cap_mim$5
Xnfet$123_0 SRLATCH_0/q vss PCP1248X$1_0/up vss nfet$123
Xnfet$123_2 SCHMITT$6_1/OUT vss fout vss nfet$123
Xnfet$123_1 SCHMITT$6_0/OUT vss foutb vss nfet$123
XNcomparator$1_0 irefn vss vdd SRLATCH_0/s Ncomparator$1_0/inn PCP1248X$1_0/out Ncomparator$1
XPcomparator$1_0 vss vdd SRLATCH_0/r irefp PCP1248X$1_0/out Pcomparator$1_0/inp Pcomparator$1
.ends

.subckt nfet$103 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$101 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt pfet$97 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$95 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt nfet$102 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$100 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt pfet$98 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$96 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt qw_NOLclk$1 VDDd VSSd PHI_2 PHI_1 CLK
Xnfet$103_1 m1_11379_n171# m1_11379_n171# VSSd VSSd m1_11837_749# VSSd nfet$103
Xnfet$103_2 m1_12351_2064# m1_12351_2064# m1_11601_2380# m1_11601_2380# m1_11837_1708#
+ VSSd nfet$103
Xnfet$103_3 m1_11161_409# m1_11161_409# VSSd VSSd m1_11837_1708# VSSd nfet$103
Xnfet$101_0 m1_12351_2064# m1_15103_233# VSSd VSSd nfet$101
Xnfet$101_1 m1_15103_233# m1_13930_233# VSSd VSSd nfet$101
Xnfet$101_2 m1_12351_431# m1_15103_1818# VSSd VSSd nfet$101
Xnfet$101_3 m1_15103_1818# m1_13930_1818# VSSd VSSd nfet$101
Xpfet$97_0 VDDd VDDd PHI_1 m1_11601_71# pfet$97
Xpfet$97_1 VDDd VDDd m1_11379_n171# m1_11161_409# pfet$97
Xpfet$97_2 VDDd VDDd PHI_2 m1_11601_2380# pfet$97
Xpfet$97_3 VDDd VDDd m1_11161_409# CLK pfet$97
Xpfet$95_0 VDDd VDDd m1_13930_233# PHI_1 pfet$95
Xpfet$95_1 VDDd VDDd m1_13930_1818# PHI_2 pfet$95
Xnfet$102_0 m1_11601_71# VSSd PHI_1 VSSd nfet$102
Xnfet$102_1 m1_11161_409# VSSd m1_11379_n171# VSSd nfet$102
Xnfet$102_2 m1_11601_2380# VSSd PHI_2 VSSd nfet$102
Xnfet$102_3 CLK VSSd m1_11161_409# VSSd nfet$102
Xnfet$100_0 PHI_1 VSSd m1_13930_233# VSSd nfet$100
Xnfet$100_1 PHI_2 VSSd m1_13930_1818# VSSd nfet$100
Xpfet$98_0 VDDd m1_11601_71# VDDd m1_11379_n171# pfet$98
Xpfet$98_1 VDDd VDDd m1_11601_71# m1_12351_431# pfet$98
Xpfet$98_2 VDDd m1_11601_2380# VDDd m1_11161_409# pfet$98
Xpfet$98_3 VDDd VDDd m1_11601_2380# m1_12351_2064# pfet$98
Xpfet$96_0 m1_12351_2064# VDDd VDDd m1_15103_233# pfet$96
Xpfet$96_1 m1_15103_233# VDDd VDDd m1_13930_233# pfet$96
Xpfet$96_2 m1_12351_431# VDDd VDDd m1_15103_1818# pfet$96
Xpfet$96_3 m1_15103_1818# VDDd VDDd m1_13930_1818# pfet$96
Xnfet$103_0 m1_12351_431# m1_12351_431# m1_11601_71# m1_11601_71# m1_11837_749# VSSd
+ nfet$103
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__latq_1$1 D E Q VDD VSS VNW VPW
X0 VSS a_1020_652# Q VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X1 a_504_110# a_36_92# VDD VNW pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X2 VDD a_1020_652# Q VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X3 a_1264_107# a_36_92# a_1020_652# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X4 VSS E a_36_92# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X5 VSS a_1364_532# a_1264_107# VPW nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X6 VDD E a_36_92# VNW pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X7 VDD a_1364_532# a_1224_652# VNW pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X8 a_872_652# D VDD VNW pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X9 a_1364_532# a_1020_652# VDD VNW pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X10 a_1020_652# a_504_110# a_872_107# VPW nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X11 a_872_107# D VSS VPW nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X12 a_1020_652# a_36_92# a_872_652# VNW pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X13 a_504_110# a_36_92# VSS VPW nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X14 a_1364_532# a_1020_652# VSS VPW nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X15 a_1224_652# a_504_110# a_1020_652# VNW pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt DFF_2phase_1$1 D Q PHI_1 PHI_2 VSSd VDDd
Xgf180mcu_fd_sc_mcu9t5v0__latq_1$1_0 gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1/Q PHI_2 Q
+ VDDd VSSd VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1$1
Xgf180mcu_fd_sc_mcu9t5v0__latq_1$1_1 D PHI_1 gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1/Q
+ VDDd VSSd VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1$1
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1$1 I VDD VSS ZN VNW VPW
X0 ZN I VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__and2_1$1 A1 A2 VDD VSS Z VNW VPW
X0 VDD A2 a_36_201# VNW pfet_05v0 ad=0.5054p pd=2.57u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1 a_244_201# A1 a_36_201# VPW nfet_05v0 ad=0.1056p pd=0.98u as=0.2904p ps=2.2u w=0.66u l=0.6u
X2 Z a_36_201# VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.3894p ps=2.06u w=1.32u l=0.6u
X3 Z a_36_201# VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.5054p ps=2.57u w=1.83u l=0.5u
X4 VSS A2 a_244_201# VPW nfet_05v0 ad=0.3894p pd=2.06u as=0.1056p ps=0.98u w=0.66u l=0.6u
X5 a_36_201# A1 VDD VNW pfet_05v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__or2_1$1 A1 A2 VDD VSS Z VNW VPW
X0 a_255_756# A1 a_67_756# VNW pfet_05v0 ad=0.2379p pd=1.435u as=0.4026p ps=2.71u w=0.915u l=0.5u
X1 VSS A2 a_67_756# VPW nfet_05v0 ad=0.3828p pd=2.08u as=0.1716p ps=1.18u w=0.66u l=0.6u
X2 VDD A2 a_255_756# VNW pfet_05v0 ad=0.57645p pd=2.69u as=0.2379p ps=1.435u w=0.915u l=0.5u
X3 Z a_67_756# VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.3828p ps=2.08u w=1.32u l=0.6u
X4 Z a_67_756# VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.57645p ps=2.69u w=1.83u l=0.5u
X5 a_67_756# A1 VSS VPW nfet_05v0 ad=0.1716p pd=1.18u as=0.2904p ps=2.2u w=0.66u l=0.6u
.ends

.subckt Register_unitcell$1 out q default phi1 en phi2 d VSSd VDDd
XDFF_2phase_1$1_0 d q phi1 phi2 VSSd VDDd DFF_2phase_1$1
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$1_0 en VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1$1
Xgf180mcu_fd_sc_mcu9t5v0__and2_1$1_0 gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN default
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1$1_0/A1 VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1$1
Xgf180mcu_fd_sc_mcu9t5v0__and2_1$1_1 q en VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1$1_0/A2
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1$1
Xgf180mcu_fd_sc_mcu9t5v0__or2_1$1_0 gf180mcu_fd_sc_mcu9t5v0__or2_1$1_0/A1 gf180mcu_fd_sc_mcu9t5v0__or2_1$1_0/A2
+ VDDd VSSd out VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1$1
.ends

.subckt SRegister_10$1 out[1] out[2] out[3] out[8] d q default10 default9 default8
+ default7 default6 default5 default4 default3 default2 default1 out[9] out[6] out[4]
+ out[10] out[7] en phi2 out[5] phi1 VSSd VDDd
XRegister_unitcell$1_0 out[2] Register_unitcell$1_7/d default2 phi1 en phi2 Register_unitcell$1_6/q
+ VSSd VDDd Register_unitcell$1
XRegister_unitcell$1_1 out[6] Register_unitcell$1_2/d default6 phi1 en phi2 Register_unitcell$1_9/q
+ VSSd VDDd Register_unitcell$1
XRegister_unitcell$1_2 out[7] Register_unitcell$1_3/d default7 phi1 en phi2 Register_unitcell$1_2/d
+ VSSd VDDd Register_unitcell$1
XRegister_unitcell$1_3 out[8] Register_unitcell$1_4/d default8 phi1 en phi2 Register_unitcell$1_3/d
+ VSSd VDDd Register_unitcell$1
XRegister_unitcell$1_4 out[9] Register_unitcell$1_5/d default9 phi1 en phi2 Register_unitcell$1_4/d
+ VSSd VDDd Register_unitcell$1
XRegister_unitcell$1_5 out[10] q default10 phi1 en phi2 Register_unitcell$1_5/d VSSd
+ VDDd Register_unitcell$1
XRegister_unitcell$1_7 out[3] Register_unitcell$1_8/d default3 phi1 en phi2 Register_unitcell$1_7/d
+ VSSd VDDd Register_unitcell$1
XRegister_unitcell$1_6 out[1] Register_unitcell$1_6/q default1 phi1 en phi2 d VSSd
+ VDDd Register_unitcell$1
XRegister_unitcell$1_8 out[4] Register_unitcell$1_9/d default4 phi1 en phi2 Register_unitcell$1_8/d
+ VSSd VDDd Register_unitcell$1
XRegister_unitcell$1_9 out[5] Register_unitcell$1_9/q default5 phi1 en phi2 Register_unitcell$1_9/d
+ VSSd VDDd Register_unitcell$1
.ends

.subckt pfet$90 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$96 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$88 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$94 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$91 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$97 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$89 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$95 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$93 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$92 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt asc_hysteresis_buffer$12 vss vdd out in
Xpfet$90_0 vdd vdd m1_348_648# in pfet$90
Xnfet$96_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$96
Xpfet$88_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd m1_884_42#
+ m1_884_42# pfet$88
Xnfet$94_0 m1_348_648# vss m1_884_42# vss nfet$94
Xpfet$91_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$91
Xnfet$97_0 m1_1156_42# vss m1_884_42# vss nfet$97
Xpfet$89_0 vdd vdd m1_884_42# m1_348_648# pfet$89
Xnfet$95_0 in vss m1_348_648# vss nfet$95
Xnfet$93_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$93
Xpfet$92_0 vdd vdd m1_884_42# m1_1156_42# pfet$92
.ends

.subckt nfet$98 a_n84_0# a_94_0# a_30_460# VSUBS
X0 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$93 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=2.6p pd=9.3u as=2.6p ps=9.3u w=4u l=0.28u
.ends

.subckt nfet$99 a_30_n132# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$94 a_28_460# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_460# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt SCHMITT$5 VDD VSS IN OUT
Xnfet$98_0 m1_592_402# OUT IN VSS nfet$98
Xnfet$98_1 VSS m1_592_402# IN VSS nfet$98
Xpfet$93_1 IN VDD VDD m1_596_1544# pfet$93
Xpfet$93_0 IN VDD m1_596_1544# OUT pfet$93
Xnfet$99_0 OUT m1_592_402# VDD VSS nfet$99
Xpfet$94_0 OUT VDD m1_596_1544# VSS pfet$94
.ends

.subckt scan_chain VDDd ENd DATAd CLKd out[1] out[2] out[3] out[4] out[5] out[6] out[7]
+ out[8] out[9] out[10] out[20] out[19] out[18] out[17] out[16] out[15] out[14] out[13]
+ out[12] out[11] out[21] out[22] out[23] out[24] out[25] out[26] out[27] out[28]
+ out[29] out[30] out[40] out[39] out[38] out[37] out[36] out[35] out[34] out[33]
+ out[32] out[31] out[41] out[42] out[43] out[44] out[45] out[46] out[47] out[48]
+ out[49] out[50] VSSd
Xqw_NOLclk$1_0 VDDd VSSd qw_NOLclk$1_0/PHI_2 qw_NOLclk$1_0/PHI_1 SCHMITT$5_0/OUT qw_NOLclk$1
XSRegister_10$1_0 out[31] out[32] out[33] out[38] SRegister_10$1_3/q SRegister_10$1_2/d
+ VSSd VSSd VDDd VSSd VSSd VDDd VDDd VSSd VSSd VSSd out[39] out[36] out[34] out[40]
+ out[37] SRegister_10$1_4/en qw_NOLclk$1_0/PHI_2 out[35] qw_NOLclk$1_0/PHI_1 VSSd
+ VDDd SRegister_10$1
XSRegister_10$1_1 out[11] out[12] out[13] out[18] SRegister_10$1_4/q SRegister_10$1_3/d
+ VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd out[19] out[16] out[14] out[20]
+ out[17] SRegister_10$1_4/en qw_NOLclk$1_0/PHI_2 out[15] qw_NOLclk$1_0/PHI_1 VSSd
+ VDDd SRegister_10$1
XSRegister_10$1_2 out[41] out[42] out[43] out[48] SRegister_10$1_2/d SRegister_10$1_2/q
+ VSSd VSSd VSSd VSSd VDDd VSSd VSSd VDDd VDDd VSSd out[49] out[46] out[44] out[50]
+ out[47] SRegister_10$1_4/en qw_NOLclk$1_0/PHI_2 out[45] qw_NOLclk$1_0/PHI_1 VSSd
+ VDDd SRegister_10$1
XSRegister_10$1_3 out[21] out[22] out[23] out[28] SRegister_10$1_3/d SRegister_10$1_3/q
+ VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd out[29] out[26] out[24] out[30]
+ out[27] SRegister_10$1_4/en qw_NOLclk$1_0/PHI_2 out[25] qw_NOLclk$1_0/PHI_1 VSSd
+ VDDd SRegister_10$1
XSRegister_10$1_4 out[1] out[2] out[3] out[8] SRegister_10$1_4/d SRegister_10$1_4/q
+ VSSd VSSd VSSd VSSd VDDd VSSd VSSd VSSd VSSd VSSd out[9] out[6] out[4] out[10] out[7]
+ SRegister_10$1_4/en qw_NOLclk$1_0/PHI_2 out[5] qw_NOLclk$1_0/PHI_1 VSSd VDDd SRegister_10$1
Xasc_hysteresis_buffer$12_0 VSSd VDDd SCHMITT$5_0/IN CLKd asc_hysteresis_buffer$12
Xasc_hysteresis_buffer$12_1 VSSd VDDd SRegister_10$1_4/en ENd asc_hysteresis_buffer$12
Xasc_hysteresis_buffer$12_2 VSSd VDDd SRegister_10$1_4/d DATAd asc_hysteresis_buffer$12
XSCHMITT$5_0 VDDd VSSd SCHMITT$5_0/IN SCHMITT$5_0/OUT SCHMITT$5
.ends

.subckt top_level_20250919_sc en clk ext_pfd_div ext_pfd_ref ext_pfd_down ext_pfd_up
+ i_cp_100u down filter_in filter_out div_in div_out ext_vco_out ext_vco_in div_def
+ up out lock data ref VSSd VDDd
Xasc_hysteresis_buffer$13_0 VSSd div_def VDDd asc_hysteresis_buffer$13_0/out asc_hysteresis_buffer$13
Xtop_level_20250912_nosc_0 i_cp_100u asc_hysteresis_buffer$13_0/out scan_chain_0/out[42]
+ scan_chain_0/out[43] scan_chain_0/out[44] scan_chain_0/out[45] scan_chain_0/out[46]
+ scan_chain_0/out[47] scan_chain_0/out[48] scan_chain_0/out[49] scan_chain_0/out[50]
+ div_out scan_chain_0/out[41] scan_chain_0/out[40] scan_chain_0/out[39] scan_chain_0/out[38]
+ scan_chain_0/out[37] scan_chain_0/out[36] scan_chain_0/out[35] scan_chain_0/out[34]
+ scan_chain_0/out[33] ref ext_pfd_div ext_pfd_ref ext_pfd_up ext_pfd_down scan_chain_0/out[1]
+ scan_chain_0/out[2] down scan_chain_0/out[6] scan_chain_0/out[5] scan_chain_0/out[4]
+ scan_chain_0/out[3] filter_in filter_out scan_chain_0/out[32] scan_chain_0/out[31]
+ scan_chain_0/out[26] scan_chain_0/out[17] scan_chain_0/out[16] scan_chain_0/out[25]
+ scan_chain_0/out[15] scan_chain_0/out[24] scan_chain_0/out[14] scan_chain_0/out[13]
+ scan_chain_0/out[12] scan_chain_0/out[11] scan_chain_0/out[10] scan_chain_0/out[9]
+ scan_chain_0/out[23] scan_chain_0/out[22] scan_chain_0/out[21] scan_chain_0/out[20]
+ scan_chain_0/out[19] scan_chain_0/out[18] scan_chain_0/out[7] scan_chain_0/out[8]
+ VCOfinal_0/fout VCOfinal_0/irefn VSSd VDDd VCOfinal_0/vin div_in ext_vco_out VCOfinal_0/irefp
+ VCOfinal_0/iref200 up lock out ext_vco_in top_level_20250912_nosc
XVCOfinal_0 VCOfinal_0/s3 VCOfinal_0/s0 VCOfinal_0/s1 VCOfinal_0/s2 VCOfinal_0/iref200
+ VCOfinal_0/fout VCOfinal_0/foutb VCOfinal_0/irefn VCOfinal_0/irefp VCOfinal_0/vin
+ VSSd VDDd VSSd VCOfinal
Xscan_chain_0 VDDd en data clk scan_chain_0/out[1] scan_chain_0/out[2] scan_chain_0/out[3]
+ scan_chain_0/out[4] scan_chain_0/out[5] scan_chain_0/out[6] scan_chain_0/out[7]
+ scan_chain_0/out[8] scan_chain_0/out[9] scan_chain_0/out[10] scan_chain_0/out[20]
+ scan_chain_0/out[19] scan_chain_0/out[18] scan_chain_0/out[17] scan_chain_0/out[16]
+ scan_chain_0/out[15] scan_chain_0/out[14] scan_chain_0/out[13] scan_chain_0/out[12]
+ scan_chain_0/out[11] scan_chain_0/out[21] scan_chain_0/out[22] scan_chain_0/out[23]
+ scan_chain_0/out[24] scan_chain_0/out[25] scan_chain_0/out[26] VCOfinal_0/s0 VCOfinal_0/s1
+ VCOfinal_0/s2 VCOfinal_0/s3 scan_chain_0/out[40] scan_chain_0/out[39] scan_chain_0/out[38]
+ scan_chain_0/out[37] scan_chain_0/out[36] scan_chain_0/out[35] scan_chain_0/out[34]
+ scan_chain_0/out[33] scan_chain_0/out[32] scan_chain_0/out[31] scan_chain_0/out[41]
+ scan_chain_0/out[42] scan_chain_0/out[43] scan_chain_0/out[44] scan_chain_0/out[45]
+ scan_chain_0/out[46] scan_chain_0/out[47] scan_chain_0/out[48] scan_chain_0/out[49]
+ scan_chain_0/out[50] VSSd scan_chain
.ends

.subckt top_level_20250919_wire ref ext_pfd_div ext_pfd_ref ext_pfd_up ext_pfd_down
+ lock i_cp_100u up down filter_in ext_vco_out ext_vco_in filter_out out div_in div_out
+ div_def clk data en VSSd VDDd
Xtop_level_20250919_sc_0 en clk ext_pfd_div ext_pfd_ref ext_pfd_down ext_pfd_up i_cp_100u
+ down filter_in filter_out div_in div_out ext_vco_out ext_vco_in div_def up out lock
+ data ref VSSd VDDd top_level_20250919_sc
.ends

