* Extracted by KLayout with GF180MCU LVS runset on : 12/08/2025 22:56

.SUBCKT xp_programmable_basic_pump VSS out down iref VDD s1 s2 s3 s4 up
M$1 VDD s1 \$37 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$2 VDD s2 \$44 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$3 VDD s3 \$38 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$4 VDD s4 \$47 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$5 VDD up \$148 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$6 \$107 \$37 \$42 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$7 iref \$37 \$66 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$8 \$107 s1 VDD VDD pfet_03v3 L=0.5U W=1U AS=0.65P AD=0.65P PS=3.3U PD=3.3U
M$9 \$108 \$44 \$42 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$10 iref \$44 \$30 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$11 \$108 s2 VDD VDD pfet_03v3 L=0.5U W=1U AS=0.65P AD=0.65P PS=3.3U PD=3.3U
M$12 \$109 \$38 \$42 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$13 iref \$38 \$4 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$14 \$109 s3 VDD VDD pfet_03v3 L=0.5U W=1U AS=0.65P AD=0.65P PS=3.3U PD=3.3U
M$15 \$147 \$47 \$42 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$16 iref \$47 \$16 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$17 \$147 s4 VDD VDD pfet_03v3 L=0.5U W=1U AS=0.65P AD=0.65P PS=3.3U PD=3.3U
M$18 VDD VDD VDD VDD pfet_03v3 L=0.5U W=252U AS=109.2P AD=109.2P PS=395.2U
+ PD=395.2U
M$19 out \$147 \$149 VDD pfet_03v3 L=0.5U W=336U AS=109.2P AD=109.2P PS=423.2U
+ PD=423.2U
M$31 out \$109 \$146 VDD pfet_03v3 L=0.5U W=168U AS=54.6P AD=54.6P PS=211.6U
+ PD=211.6U
M$57 \$149 \$148 VDD VDD pfet_03v3 L=0.5U W=336U AS=109.2P AD=109.2P PS=423.2U
+ PD=423.2U
M$69 \$146 \$148 VDD VDD pfet_03v3 L=0.5U W=168U AS=54.6P AD=54.6P PS=211.6U
+ PD=211.6U
M$101 \$168 \$148 VDD VDD pfet_03v3 L=0.5U W=84U AS=27.3P AD=27.3P PS=105.8U
+ PD=105.8U
M$107 \$170 \$148 VDD VDD pfet_03v3 L=0.5U W=42U AS=13.65P AD=13.65P PS=52.9U
+ PD=52.9U
M$113 \$169 VSS VDD VDD pfet_03v3 L=0.5U W=42U AS=13.65P AD=13.65P PS=52.9U
+ PD=52.9U
M$139 out \$108 \$168 VDD pfet_03v3 L=0.5U W=84U AS=27.3P AD=27.3P PS=105.8U
+ PD=105.8U
M$145 out \$107 \$170 VDD pfet_03v3 L=0.5U W=42U AS=13.65P AD=13.65P PS=52.9U
+ PD=52.9U
M$151 \$42 \$42 \$169 VDD pfet_03v3 L=0.5U W=42U AS=13.65P AD=13.65P PS=52.9U
+ PD=52.9U
M$246 VSS VSS VSS VSS nfet_03v3 L=0.5U W=168U AS=73.08P AD=73.08P PS=272.88U
+ PD=272.88U
M$248 out \$16 \$17 VSS nfet_03v3 L=0.5U W=112U AS=48.72P AD=48.72P PS=181.92U
+ PD=181.92U
M$252 out \$4 \$5 VSS nfet_03v3 L=0.5U W=56U AS=24.36P AD=24.36P PS=90.96U
+ PD=90.96U
M$264 \$17 down VSS VSS nfet_03v3 L=0.5U W=112U AS=48.72P AD=48.72P PS=181.92U
+ PD=181.92U
M$268 \$5 down VSS VSS nfet_03v3 L=0.5U W=56U AS=24.36P AD=24.36P PS=90.96U
+ PD=90.96U
M$280 \$29 down VSS VSS nfet_03v3 L=0.5U W=28U AS=12.18P AD=12.18P PS=45.48U
+ PD=45.48U
M$282 \$39 VDD VSS VSS nfet_03v3 L=0.5U W=14U AS=6.09P AD=6.09P PS=22.74U
+ PD=22.74U
M$284 \$40 down VSS VSS nfet_03v3 L=0.5U W=14U AS=6.09P AD=6.09P PS=22.74U
+ PD=22.74U
M$286 \$41 VDD VSS VSS nfet_03v3 L=0.5U W=14U AS=6.09P AD=6.09P PS=22.74U
+ PD=22.74U
M$294 out \$30 \$29 VSS nfet_03v3 L=0.5U W=28U AS=12.18P AD=12.18P PS=45.48U
+ PD=45.48U
M$296 iref iref \$39 VSS nfet_03v3 L=0.5U W=14U AS=6.09P AD=6.09P PS=22.74U
+ PD=22.74U
M$298 out \$66 \$40 VSS nfet_03v3 L=0.5U W=14U AS=6.09P AD=6.09P PS=22.74U
+ PD=22.74U
M$300 \$42 iref \$41 VSS nfet_03v3 L=0.5U W=14U AS=6.09P AD=6.09P PS=22.74U
+ PD=22.74U
M$322 VSS \$37 \$66 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$323 iref s1 \$66 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$324 VSS s1 \$37 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$325 VSS \$44 \$30 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$326 iref s2 \$30 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$327 VSS s2 \$44 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$328 VSS \$38 \$4 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$329 VSS s3 \$38 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$330 iref s3 \$4 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$331 VSS \$47 \$16 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$332 VSS s4 \$47 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$333 iref s4 \$16 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$334 VSS up \$148 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$351 \$107 s1 \$42 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$352 \$108 s2 \$42 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$353 \$109 s3 \$42 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$354 \$147 s4 \$42 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
.ENDS xp_programmable_basic_pump
