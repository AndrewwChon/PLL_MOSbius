* Extracted by KLayout with GF180MCU LVS runset on : 07/08/2025 03:02

.SUBCKT asc_NOR VSS A OUT B VDD
M$1 \$10 A VDD VDD pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U PD=13.3U
M$2 OUT B \$10 VDD pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U PD=13.3U
M$3 OUT A VSS VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$4 VSS B OUT VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
.ENDS asc_NOR
