* NGSPICE file created from xp_programmable_basic_pump.ext - technology: gf180mcuD

.subckt nfet$2 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$3 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_954_0# w_n180_n88# a_854_n136#
+ a_n92_0# a_446_n136# a_650_n136# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt nfet$1$1 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$6 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$4 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt inv1u05u VDD in VSS out
Xpfet$6_0 VDD VDD out in pfet$6
Xnfet$4_0 in VSS out VSS nfet$4
.ends

.subckt pfet$4 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.5u
.ends

.subckt pfet$7 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$6 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pass1u05u VDD VSS ind ins clkp clkn
Xpfet$7_0 VDD ind ins clkp pfet$7
Xnfet$6_0 clkn ind ins VSS nfet$6
.ends

.subckt pfet$2 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=4.55p ps=15.3u w=7u l=0.5u
.ends

.subckt nfet$5 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$1$1 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_954_0# w_n180_n88#
+ a_38_n60# a_n92_0# a_1058_n60# a_854_n60# a_342_0# a_138_0# a_650_n60#
X0 a_954_0# a_854_n60# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n60# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt nfet$2$1 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt xp_programmable_basic_pump up vss vdd s1 s2 s3 s4 down out iref
Xnfet$2_2 vss down vss m1_n7879_n12170# down vss nfet$2
Xpfet$3_9 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$3
Xnfet$2_15 vss down vss m1_n8607_n8040# down vss nfet$2
Xnfet$1$1_1 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$1$1
Xinv1u05u_3 vdd s1 vss inv1u05u_3/out inv1u05u
Xnfet$2_3 vss down vss m1_n7879_n12170# down vss nfet$2
Xnfet$1$1_2 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$1$1
Xnfet$2_4 vss down vss m1_n7879_n12170# down vss nfet$2
Xnfet$1$1_10 pass1u05u_2/ins pass1u05u_2/ins m1_n7679_n8960# m1_n7679_n8960# out vss
+ nfet$1$1
Xnfet$1$1_3 vss vss vss vss vss vss nfet$1$1
Xnfet$2_5 vss down vss m1_n7879_n12170# down vss nfet$2
Xnfet$1$1_11 vss vss vss vss vss vss nfet$1$1
Xnfet$1$1_4 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$1$1
Xnfet$2_6 m1_n7879_n12170# pass1u05u_0/ins m1_n7879_n12170# out pass1u05u_0/ins vss
+ nfet$2
Xnfet$1$1_12 down down vss vss m1_n7679_n8960# vss nfet$1$1
Xnfet$1$1_5 vss vss vss vss vss vss nfet$1$1
Xnfet$2_7 m1_n7879_n12170# pass1u05u_0/ins m1_n7879_n12170# out pass1u05u_0/ins vss
+ nfet$2
Xnfet$1$1_13 vss vss vss vss vss vss nfet$1$1
Xnfet$1$1_6 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$1$1
Xnfet$2_8 vss vdd vss m1_n8144_n9165# vdd vss nfet$2
Xnfet$1$1_14 vss vss vss vss vss vss nfet$1$1
Xnfet$1$1_7 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$1$1
Xnfet$2_9 m1_n7216_n8262# iref m1_n7216_n8262# pass1u05u_7/ind iref vss nfet$2
Xnfet$1$1_15 vss vss vss vss vss vss nfet$1$1
Xnfet$1$1_8 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$1$1
Xpfet$4_0 vdd s3 pass1u05u_5/ins vdd pfet$4
Xnfet$1$1_9 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$1$1
Xpfet$4_1 vdd s2 pass1u05u_4/ins vdd pfet$4
Xpfet$4_2 vdd s1 pass1u05u_3/ins vdd pfet$4
Xpfet$4_3 vdd s4 pass1u05u_7/ins vdd pfet$4
Xpass1u05u_0 vdd vss iref pass1u05u_0/ins inv1u05u_1/out s3 pass1u05u
Xpfet$2_0 vdd vdd vdd vdd pfet$2
Xnfet$5_0 inv1u05u_2/out pass1u05u_1/ins vss vss nfet$5
Xpfet$2_20 vdd vdd vdd vdd pfet$2
Xpass1u05u_1 vdd vss iref pass1u05u_1/ins inv1u05u_2/out s2 pass1u05u
Xpfet$2_1 vdd vdd vdd vdd pfet$2
Xnfet$5_1 inv1u05u_3/out pass1u05u_2/ins vss vss nfet$5
Xpfet$2_2 vdd vdd vdd vdd pfet$2
Xpfet$2_21 vdd vdd vdd vdd pfet$2
Xpass1u05u_2 vdd vss iref pass1u05u_2/ins inv1u05u_3/out s1 pass1u05u
Xpfet$2_10 vdd vdd vdd vdd pfet$2
Xnfet$5_2 inv1u05u_0/out pass1u05u_6/ins vss vss nfet$5
Xpfet$2_3 vdd vdd vdd vdd pfet$2
Xpfet$2_11 vdd vdd vdd vdd pfet$2
Xpfet$2_22 vdd vdd vdd vdd pfet$2
Xpass1u05u_3 vdd vss pass1u05u_7/ind pass1u05u_3/ins inv1u05u_3/out s1 pass1u05u
Xpfet$1$1_0 vdd vdd m1_n4127_3649# vss vss m1_n4127_3649# vdd vss vdd vss vss vdd
+ m1_n4127_3649# vss pfet$1$1
Xnfet$5_3 inv1u05u_1/out pass1u05u_0/ins vss vss nfet$5
Xpass1u05u_4 vdd vss pass1u05u_7/ind pass1u05u_4/ins inv1u05u_2/out s2 pass1u05u
Xpfet$2_12 vdd vdd vdd vdd pfet$2
Xpfet$2_4 vdd vdd vdd vdd pfet$2
Xpfet$2_23 vdd vdd vdd vdd pfet$2
Xpfet$1$1_1 m1_n5580_883# m1_n5580_883# out pass1u05u_5/ins pass1u05u_5/ins out vdd
+ pass1u05u_5/ins m1_n5580_883# pass1u05u_5/ins pass1u05u_5/ins m1_n5580_883# out
+ pass1u05u_5/ins pfet$1$1
Xpfet$2_13 vdd vdd vdd vdd pfet$2
Xpass1u05u_5 vdd vss pass1u05u_7/ind pass1u05u_5/ins inv1u05u_1/out s3 pass1u05u
Xpfet$2_5 vdd vdd vdd vdd pfet$2
Xpfet$1$1_2 m1_n5580_883# m1_n5580_883# out pass1u05u_5/ins pass1u05u_5/ins out vdd
+ pass1u05u_5/ins m1_n5580_883# pass1u05u_5/ins pass1u05u_5/ins m1_n5580_883# out
+ pass1u05u_5/ins pfet$1$1
Xpfet$2_14 vdd vdd vdd vdd pfet$2
Xpass1u05u_6 vdd vss iref pass1u05u_6/ins inv1u05u_0/out s4 pass1u05u
Xpfet$2_6 vdd vdd vdd vdd pfet$2
Xpfet$1$1_3 m1_n5580_883# m1_n5580_883# out pass1u05u_5/ins pass1u05u_5/ins out vdd
+ pass1u05u_5/ins m1_n5580_883# pass1u05u_5/ins pass1u05u_5/ins m1_n5580_883# out
+ pass1u05u_5/ins pfet$1$1
Xpfet$2_15 vdd vdd vdd vdd pfet$2
Xpass1u05u_7 vdd vss pass1u05u_7/ind pass1u05u_7/ins inv1u05u_0/out s4 pass1u05u
Xpfet$2_7 vdd vdd vdd vdd pfet$2
Xpfet$1$1_4 m1_n5580_883# m1_n5580_883# out pass1u05u_5/ins pass1u05u_5/ins out vdd
+ pass1u05u_5/ins m1_n5580_883# pass1u05u_5/ins pass1u05u_5/ins m1_n5580_883# out
+ pass1u05u_5/ins pfet$1$1
Xpfet$2_16 vdd vdd vdd vdd pfet$2
Xpfet$2_8 vdd vdd vdd vdd pfet$2
Xpfet$1$1_5 m1_n4127_3649# m1_n4127_3649# pass1u05u_7/ind pass1u05u_7/ind pass1u05u_7/ind
+ pass1u05u_7/ind vdd pass1u05u_7/ind m1_n4127_3649# pass1u05u_7/ind pass1u05u_7/ind
+ m1_n4127_3649# pass1u05u_7/ind pass1u05u_7/ind pfet$1$1
Xpfet$2_17 vdd vdd vdd vdd pfet$2
Xpfet$2_9 vdd vdd vdd vdd pfet$2
Xpfet$2_18 vdd vdd vdd vdd pfet$2
Xpfet$2_19 vdd vdd vdd vdd pfet$2
Xpfet$3_20 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$3
Xnfet$2$1_0 down down vss vss m1_n8807_n11192# vss nfet$2$1
Xpfet$3_10 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$3
Xpfet$3_21 m1_n6703_2564# m1_n6703_2564# pass1u05u_4/ins out out vdd pass1u05u_4/ins
+ m1_n6703_2564# pass1u05u_4/ins pass1u05u_4/ins m1_n6703_2564# out pass1u05u_4/ins
+ pass1u05u_4/ins pfet$3
Xnfet$2$1_1 down down vss vss m1_n8807_n11192# vss nfet$2$1
Xpfet$3_22 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$3
Xpfet$3_11 vdd vdd up m1_n5450_4559# m1_n5450_4559# vdd up vdd up up vdd m1_n5450_4559#
+ up up pfet$3
Xnfet$2$1_2 down down vss vss m1_n8807_n11192# vss nfet$2$1
Xpfet$3_23 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$3
Xpfet$3_12 vdd vdd up m1_n6703_2564# m1_n6703_2564# vdd up vdd up up vdd m1_n6703_2564#
+ up up pfet$3
Xnfet$2$1_10 vss vss vss vss vss vss nfet$2$1
Xpfet$3_0 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$3
Xnfet$2$1_3 down down vss vss m1_n8807_n11192# vss nfet$2$1
Xpfet$3_24 m1_n5450_4559# m1_n5450_4559# pass1u05u_3/ins out out vdd pass1u05u_3/ins
+ m1_n5450_4559# pass1u05u_3/ins pass1u05u_3/ins m1_n5450_4559# out pass1u05u_3/ins
+ pass1u05u_3/ins pfet$3
Xpfet$3_13 vdd vdd up m1_n6703_2564# m1_n6703_2564# vdd up vdd up up vdd m1_n6703_2564#
+ up up pfet$3
Xnfet$2$1_11 vss vss vss vss vss vss nfet$2$1
Xpfet$3_1 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$3
Xnfet$2$1_4 vss vss vss vss vss vss nfet$2$1
Xpfet$3_25 m1_n6703_2564# m1_n6703_2564# pass1u05u_4/ins out out vdd pass1u05u_4/ins
+ m1_n6703_2564# pass1u05u_4/ins pass1u05u_4/ins m1_n6703_2564# out pass1u05u_4/ins
+ pass1u05u_4/ins pfet$3
Xpfet$3_14 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$3
Xnfet$2$1_12 vss vss vss vss vss vss nfet$2$1
Xpfet$3_2 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$3
Xnfet$2$1_5 vss vss vss vss vss vss nfet$2$1
Xpfet$3_15 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$3
Xnfet$2$1_13 vss vss vss vss vss vss nfet$2$1
Xpfet$3_3 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$3
Xnfet$2$1_6 down down vss vss m1_n8807_n11192# vss nfet$2$1
Xpfet$3_16 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$3
Xnfet$2_10 m1_n8607_n8040# pass1u05u_1/ins m1_n8607_n8040# out pass1u05u_1/ins vss
+ nfet$2
Xpfet$3_4 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$3
Xnfet$2$1_7 down down vss vss m1_n8807_n11192# vss nfet$2$1
Xpfet$3_17 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$3
Xpfet$3_5 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$3
Xnfet$2_11 m1_n8144_n9165# iref m1_n8144_n9165# iref iref vss nfet$2
Xnfet$2$1_8 down down vss vss m1_n8807_n11192# vss nfet$2$1
Xpfet$3_18 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$3
Xpfet$3_6 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$3
Xnfet$2_12 vss down vss m1_n8607_n8040# down vss nfet$2
Xinv1u05u_0 vdd s4 vss inv1u05u_0/out inv1u05u
Xnfet$2$1_9 down down vss vss m1_n8807_n11192# vss nfet$2$1
Xpfet$3_19 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$3
Xnfet$2_0 m1_n7879_n12170# pass1u05u_0/ins m1_n7879_n12170# out pass1u05u_0/ins vss
+ nfet$2
Xpfet$3_7 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$3
Xnfet$2_13 vss vdd vss m1_n7216_n8262# vdd vss nfet$2
Xinv1u05u_1 vdd s3 vss inv1u05u_1/out inv1u05u
Xpfet$3_8 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$3
Xnfet$2_1 m1_n7879_n12170# pass1u05u_0/ins m1_n7879_n12170# out pass1u05u_0/ins vss
+ nfet$2
Xnfet$2_14 m1_n8607_n8040# pass1u05u_1/ins m1_n8607_n8040# out pass1u05u_1/ins vss
+ nfet$2
Xnfet$1$1_0 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out
+ vss nfet$1$1
Xinv1u05u_2 vdd s2 vss inv1u05u_2/out inv1u05u
.ends

