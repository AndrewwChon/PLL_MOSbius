** sch_path: /foss/designs/libs/secondary_esd/io_secondary_3p3.sch
.subckt io_secondary_3p3 VDD to_gate ASIG3V3 VSS
*.PININFO VSS:B VDD:B to_gate:B ASIG3V3:B
XR1 to_gate ASIG3V3 VSS ppolyf_u r_width=40e-6 r_length=5.5e-6 m=1
D2 VSS to_gate diode_nd2ps_03v3 area='10u * 10u ' pj='2*10u + 2*10u ' m=4
D1 to_gate VDD diode_pd2nw_03v3 area='10u * 10u ' pj='2*10u + 2*10u ' m=4
.ends
