* NGSPICE file created from top_level_20250919_final.ext - technology: gf180mcuD

.subckt ppolyf_u_resistor$6 a_n376_0# a_5400_0# a_n132_0#
X0 a_n132_0# a_5400_0# a_n376_0# ppolyf_u r_width=1u r_length=27u
.ends

.subckt cap_nmos a_88_n92# a_0_0#
X0 a_88_n92# a_0_0# cap_nmos_03v3 c_width=10u c_length=10u
.ends

.subckt DECAP_SC a_n313_2257# vdd vss
Xcap_nmos_0 vdd vss cap_nmos
Xcap_nmos_1 vdd vss cap_nmos
Xcap_nmos_2 vdd vss cap_nmos
Xcap_nmos_3 vdd vss cap_nmos
.ends

.subckt DECAP_LARGE vdd vss
XDECAP_SC_0 vss vdd vss DECAP_SC
XDECAP_SC_1 vss vdd vss DECAP_SC
XDECAP_SC_2 DECAP_SC_2/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_3 DECAP_SC_3/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_4 DECAP_SC_4/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_5 DECAP_SC_5/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_6 DECAP_SC_6/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_7 DECAP_SC_7/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_8 DECAP_SC_8/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_90 DECAP_SC_90/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_9 DECAP_SC_9/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_80 vss vdd vss DECAP_SC
XDECAP_SC_91 DECAP_SC_91/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_70 vss vdd vss DECAP_SC
XDECAP_SC_81 vss vdd vss DECAP_SC
XDECAP_SC_92 vss vdd vss DECAP_SC
XDECAP_SC_71 vss vdd vss DECAP_SC
XDECAP_SC_60 vss vdd vss DECAP_SC
XDECAP_SC_93 vss vdd vss DECAP_SC
XDECAP_SC_82 vss vdd vss DECAP_SC
XDECAP_SC_50 vss vdd vss DECAP_SC
XDECAP_SC_72 DECAP_SC_72/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_94 vss vdd vss DECAP_SC
XDECAP_SC_61 vss vdd vss DECAP_SC
XDECAP_SC_83 vss vdd vss DECAP_SC
XDECAP_SC_40 DECAP_SC_40/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_51 vss vdd vss DECAP_SC
XDECAP_SC_73 vss vdd vss DECAP_SC
XDECAP_SC_95 vss vdd vss DECAP_SC
XDECAP_SC_62 vss vdd vss DECAP_SC
XDECAP_SC_84 vss vdd vss DECAP_SC
XDECAP_SC_52 DECAP_SC_52/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_41 DECAP_SC_41/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_30 vss vdd vss DECAP_SC
XDECAP_SC_120 DECAP_SC_120/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_96 DECAP_SC_96/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_63 vss vdd vss DECAP_SC
XDECAP_SC_74 vss vdd vss DECAP_SC
XDECAP_SC_85 vss vdd vss DECAP_SC
XDECAP_SC_64 vss vdd vss DECAP_SC
XDECAP_SC_42 vss vdd vss DECAP_SC
XDECAP_SC_31 vss vdd vss DECAP_SC
XDECAP_SC_20 vss vdd vss DECAP_SC
XDECAP_SC_97 vss vdd vss DECAP_SC
XDECAP_SC_53 vss vdd vss DECAP_SC
XDECAP_SC_75 vss vdd vss DECAP_SC
XDECAP_SC_86 vss vdd vss DECAP_SC
XDECAP_SC_121 vss vdd vss DECAP_SC
XDECAP_SC_110 vss vdd vss DECAP_SC
XDECAP_SC_65 vss vdd vss DECAP_SC
XDECAP_SC_43 vss vdd vss DECAP_SC
XDECAP_SC_54 vss vdd vss DECAP_SC
XDECAP_SC_21 vss vdd vss DECAP_SC
XDECAP_SC_10 vss vdd vss DECAP_SC
XDECAP_SC_122 vss vdd vss DECAP_SC
XDECAP_SC_98 vss vdd vss DECAP_SC
XDECAP_SC_100 vss vdd vss DECAP_SC
XDECAP_SC_111 vss vdd vss DECAP_SC
XDECAP_SC_32 DECAP_SC_32/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_76 vss vdd vss DECAP_SC
XDECAP_SC_87 vss vdd vss DECAP_SC
XDECAP_SC_66 vss vdd vss DECAP_SC
XDECAP_SC_44 DECAP_SC_44/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_88 vss vdd vss DECAP_SC
XDECAP_SC_55 vss vdd vss DECAP_SC
XDECAP_SC_22 vss vdd vss DECAP_SC
XDECAP_SC_11 vss vdd vss DECAP_SC
XDECAP_SC_99 vss vdd vss DECAP_SC
XDECAP_SC_33 vss vdd vss DECAP_SC
XDECAP_SC_77 vss vdd vss DECAP_SC
XDECAP_SC_123 vss vdd vss DECAP_SC
XDECAP_SC_101 vss vdd vss DECAP_SC
XDECAP_SC_112 DECAP_SC_112/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_67 vss vdd vss DECAP_SC
XDECAP_SC_89 vss vdd vss DECAP_SC
XDECAP_SC_56 vss vdd vss DECAP_SC
XDECAP_SC_23 vss vdd vss DECAP_SC
XDECAP_SC_12 DECAP_SC_12/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_102 DECAP_SC_102/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_124 vss vdd vss DECAP_SC
XDECAP_SC_113 vss vdd vss DECAP_SC
XDECAP_SC_34 vss vdd vss DECAP_SC
XDECAP_SC_45 DECAP_SC_45/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_78 vss vdd vss DECAP_SC
XDECAP_SC_46 vss vdd vss DECAP_SC
XDECAP_SC_68 vss vdd vss DECAP_SC
XDECAP_SC_57 vss vdd vss DECAP_SC
XDECAP_SC_24 vss vdd vss DECAP_SC
XDECAP_SC_13 vss vdd vss DECAP_SC
XDECAP_SC_103 DECAP_SC_103/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_125 vss vdd vss DECAP_SC
XDECAP_SC_114 vss vdd vss DECAP_SC
XDECAP_SC_35 vss vdd vss DECAP_SC
XDECAP_SC_79 vss vdd vss DECAP_SC
XDECAP_SC_47 vss vdd vss DECAP_SC
XDECAP_SC_69 vss vdd vss DECAP_SC
XDECAP_SC_25 vss vdd vss DECAP_SC
XDECAP_SC_14 vss vdd vss DECAP_SC
XDECAP_SC_58 vss vdd vss DECAP_SC
XDECAP_SC_36 vss vdd vss DECAP_SC
XDECAP_SC_104 DECAP_SC_104/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_115 vss vdd vss DECAP_SC
XDECAP_SC_48 vss vdd vss DECAP_SC
XDECAP_SC_26 vss vdd vss DECAP_SC
XDECAP_SC_15 vss vdd vss DECAP_SC
XDECAP_SC_105 DECAP_SC_105/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_116 vss vdd vss DECAP_SC
XDECAP_SC_59 DECAP_SC_59/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_37 vss vdd vss DECAP_SC
XDECAP_SC_49 vss vdd vss DECAP_SC
XDECAP_SC_27 vss vdd vss DECAP_SC
XDECAP_SC_16 vss vdd vss DECAP_SC
XDECAP_SC_38 vss vdd vss DECAP_SC
XDECAP_SC_106 DECAP_SC_106/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_117 vss vdd vss DECAP_SC
XDECAP_SC_28 vss vdd vss DECAP_SC
XDECAP_SC_17 vss vdd vss DECAP_SC
XDECAP_SC_107 DECAP_SC_107/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_118 vss vdd vss DECAP_SC
XDECAP_SC_39 vss vdd vss DECAP_SC
XDECAP_SC_29 vss vdd vss DECAP_SC
XDECAP_SC_18 vss vdd vss DECAP_SC
XDECAP_SC_108 DECAP_SC_108/a_n313_2257# vdd vss DECAP_SC
XDECAP_SC_119 vss vdd vss DECAP_SC
XDECAP_SC_19 vss vdd vss DECAP_SC
XDECAP_SC_109 DECAP_SC_109/a_n313_2257# vdd vss DECAP_SC
.ends

.subckt diode_nd2ps a_n168_0# a_0_0#
D0 a_n168_0# a_0_0# diode_nd2ps_03v3 pj=40u area=99.99999p
.ends

.subckt diode_pd2nw w_n224_n86# a_0_0#
D0 a_0_0# w_n224_n86# diode_pd2nw_03v3 pj=40u area=99.99999p
.ends

.subckt ppolyf_u_resistor$3 a_n376_0# a_1100_0# a_n132_0#
X0 a_n132_0# a_1100_0# a_n376_0# ppolyf_u r_width=40u r_length=5.5u
.ends

.subckt io_secondary_3p3 ASIG3V3 VDD VSS to_gate
Xdiode_nd2ps_0 VSS to_gate diode_nd2ps
Xdiode_nd2ps_1 VSS to_gate diode_nd2ps
Xdiode_pd2nw_0 VDD to_gate diode_pd2nw
Xdiode_nd2ps_2 VSS to_gate diode_nd2ps
Xdiode_pd2nw_1 VDD to_gate diode_pd2nw
Xdiode_nd2ps_3 VSS to_gate diode_nd2ps
Xdiode_pd2nw_2 VDD to_gate diode_pd2nw
Xdiode_pd2nw_3 VDD to_gate diode_pd2nw
Xppolyf_u_resistor$3_0 VSS ASIG3V3 to_gate ppolyf_u_resistor$3
.ends

.subckt pfet$270 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$287 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$285 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$268 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$266 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$288 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$286 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$284 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$269 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$267 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt asc_hysteresis_buffer$4 vss in vdd out
Xpfet$270_0 vdd vdd m1_884_42# m1_1156_42# pfet$270
Xnfet$287_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$287
Xnfet$285_0 m1_348_648# vss m1_884_42# vss nfet$285
Xpfet$268_0 vdd vdd m1_348_648# in pfet$268
Xpfet$266_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd
+ m1_884_42# m1_884_42# pfet$266
Xnfet$288_0 m1_1156_42# vss m1_884_42# vss nfet$288
Xnfet$286_0 in vss m1_348_648# vss nfet$286
Xnfet$284_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$284
Xpfet$269_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$269
Xpfet$267_0 vdd vdd m1_884_42# m1_348_648# pfet$267
.ends

.subckt pfet$286 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$305 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$287 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$304 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt xp_3_1_MUX$3 S0 S1 VDD VSS OUT_1 C_1 B_1 A_1
Xpfet$286_0 VDD A_1 m1_239_n318# m1_n432_458# pfet$286
Xpfet$286_2 VDD B_1 m1_239_n318# S0 pfet$286
Xpfet$286_1 VDD C_1 OUT_1 S1 pfet$286
Xpfet$286_3 VDD m1_239_n318# OUT_1 m1_n432_n1290# pfet$286
Xnfet$305_0 S1 VSS m1_n432_n1290# VSS nfet$305
Xnfet$305_1 S0 VSS m1_n432_458# VSS nfet$305
Xpfet$287_0 VDD VDD m1_n432_n1290# S1 pfet$287
Xpfet$287_1 VDD VDD m1_n432_458# S0 pfet$287
Xnfet$304_0 m1_n432_n1290# C_1 OUT_1 VSS nfet$304
Xnfet$304_1 m1_n432_458# B_1 m1_239_n318# VSS nfet$304
Xnfet$304_2 S1 m1_239_n318# OUT_1 VSS nfet$304
Xnfet$304_3 S0 A_1 m1_239_n318# VSS nfet$304
.ends

.subckt nfet$242 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$245 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$251 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$228 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$247 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$250 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$242 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$235 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$244 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$269 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$232 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$227 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$249 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$268 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$241 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$254 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$261 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$239 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$253 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$243 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$273 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$258 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$240 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$266 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$233 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$259 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$256 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$271 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$264 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$249 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$231 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$257 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$254 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$262 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$247 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$230 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$255 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$248 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$252 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$260 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$245 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$238 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$253 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$246 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$250 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$276 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$243 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$251 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$236 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$229 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$259 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$274 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$241 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$267 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$234 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$272 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$257 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$265 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$258 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$270 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$255 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$263 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$248 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$256 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$246 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$277 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$244 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$252 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$237 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$275 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_dual_psd_def_20250809$3 vdd vss pd1 pd2 pd3 pd4 pd5 pd6 pd7 pd8 pd9 fout
+ sd1 sd2 sd3 sd4 sd5 sd6 sd7 sd8 sd9 fin define
Xnfet$242_80 m1_28147_25662# m1_28991_24224# m1_30095_25658# vss nfet$242
Xnfet$245_2 m1_6275_17836# m1_7555_16080# m1_7088_18030# vss nfet$245
Xpfet$251_5 vdd vdd m1_n10308_24542# m1_n9952_24224# pfet$251
Xpfet$228_109 vdd vdd m1_10299_17343# m1_13198_17714# pfet$228
Xnfet$247_14 m1_21564_17714# vss m1_23486_19550# vss nfet$247
Xnfet$250_0 m1_n10452_25858# vss m1_n1271_25858# vss nfet$250
Xpfet$242_1 vdd m1_35837_22102# m1_35837_22102# m1_36073_22344# fout fout pfet$242
Xpfet$235_0 vdd vdd m1_n647_25662# m1_n789_25858# pfet$235
Xnfet$244_15 m1_21564_17714# m1_21564_17714# vss vss m1_24556_20470# vss nfet$244
Xnfet$269_12 m1_n10452_25858# vss m1_n5571_25662# vss nfet$269
Xpfet$232_10 vdd vdd m1_27031_17343# m1_n10452_25858# pfet$232
Xpfet$227_65 vdd vdd m1_18073_21786# m1_20126_25858# pfet$227
Xpfet$227_54 vdd vdd m1_24808_24224# m1_24188_23922# pfet$227
Xpfet$227_43 vdd vdd m1_12805_21786# pd5 pfet$227
Xnfet$245_80 m1_18824_17836# m1_19747_15778# m1_18926_16202# vss nfet$245
Xnfet$249_9 m1_n10452_25858# vss m1_27031_17343# vss nfet$249
Xpfet$227_32 vdd vdd m1_7720_24542# m1_8076_24224# pfet$227
Xpfet$227_21 vdd m1_7456_23922# m1_7720_24542# m1_7095_25858# pfet$227
Xpfet$227_10 vdd m1_8076_24224# m1_9180_25658# m1_7095_25858# pfet$227
Xnfet$268_1 m1_n1927_20274# m1_n1927_20274# vss vss m1_n2445_20470# vss nfet$268
Xnfet$241_27 m1_12875_24346# m1_12875_24346# vss vss m1_12357_24542# vss nfet$241
Xpfet$227_98 vdd m1_30095_25658# m1_30888_24542# m1_28147_25662# pfet$227
Xpfet$227_87 vdd vdd m1_28147_25662# m1_28010_25858# pfet$227
Xpfet$227_76 vdd m1_20005_23922# m1_20269_24542# m1_19644_25858# pfet$227
Xnfet$241_16 m1_24808_24224# m1_24808_24224# m1_24452_24542# m1_24452_24542# m1_24906_24542#
+ vss nfet$241
Xnfet$254_7 m1_488_21786# m1_488_21786# vss vss m1_n674_21586# vss nfet$254
Xnfet$247_6 m1_9015_17714# vss m1_12935_19550# vss nfet$247
Xnfet$261_8 m1_3015_15778# m1_3015_15778# m1_2905_18030# m1_2905_18030# m1_3141_17358#
+ vss nfet$261
Xpfet$239_7 vdd m1_32554_23922# m1_32818_24542# m1_32193_25858# pfet$239
Xpfet$253_9 vdd vdd m1_n4464_25980# m1_n4623_25487# pfet$253
Xnfet$242_81 m1_n7513_20152# vss m1_25424_24346# vss nfet$242
Xnfet$242_70 m1_21590_21786# vss m1_28010_25858# vss nfet$242
Xnfet$245_3 m1_n7513_20152# vss m1_9944_16080# vss nfet$245
Xnfet$247_15 m1_17697_15478# vss m1_22205_20152# vss nfet$247
Xpfet$251_6 vdd m1_n10308_24542# vdd m1_n9336_24346# pfet$251
Xpfet$227_110 vdd m1_11903_24542# vdd m1_12875_24346# pfet$227
Xpfet$235_10 vdd vdd m1_35071_24542# m1_32675_25947# pfet$235
Xnfet$243_0 m1_n1133_21590# m1_n1133_21590# m1_354_22513# m1_354_22513# m1_n674_21586#
+ vss nfet$243
Xpfet$235_1 vdd vdd m1_n1134_25662# m1_n1271_25858# pfet$235
Xnfet$250_1 m1_n789_25858# vss m1_n647_25662# vss nfet$250
Xpfet$228_0 vdd vdd m1_12355_15778# m1_9485_17714# pfet$228
Xnfet$244_16 m1_23486_19550# m1_23486_19550# vss vss m1_23924_20470# vss nfet$244
Xnfet$269_13 fin vss m1_n4623_25487# vss nfet$269
Xpfet$232_11 vdd vdd m1_26807_17518# m1_26217_17714# pfet$232
Xnfet$245_81 m1_13198_17714# vss m1_10299_17343# vss nfet$245
Xnfet$245_70 m1_n7513_20152# vss m1_18310_16080# vss nfet$245
Xpfet$227_99 vdd vdd m1_26705_24542# m1_24309_25858# pfet$227
Xpfet$227_88 vdd vdd m1_28634_25662# m1_28492_25858# pfet$227
Xpfet$227_77 vdd vdd m1_20269_24542# m1_20625_24224# pfet$227
Xpfet$227_66 vdd vdd m1_15461_25858# m1_11039_21786# pfet$227
Xpfet$227_55 vdd m1_24451_25662# m1_24188_23922# m1_23964_25662# pfet$227
Xnfet$241_17 m1_20625_24224# m1_20625_24224# m1_20269_24542# m1_20269_24542# m1_20723_24542#
+ vss nfet$241
Xpfet$227_44 vdd m1_15943_25858# vdd m1_17546_25658# pfet$227
Xpfet$227_33 vdd vdd m1_7522_21786# m1_7577_25858# pfet$227
Xpfet$227_22 vdd vdd m1_3537_24542# m1_3893_24224# pfet$227
Xpfet$227_11 vdd vdd m1_7719_25662# m1_7577_25858# pfet$227
Xnfet$268_2 m1_n3206_20274# m1_n3206_20274# vss vss m1_n3724_20470# vss nfet$268
Xnfet$261_9 m1_2194_16202# m1_2194_16202# vss vss m1_1676_16398# vss nfet$261
Xnfet$254_8 m1_25739_21786# m1_25739_21786# vss vss m1_24577_21586# vss nfet$254
Xnfet$247_7 m1_5148_15478# vss m1_11654_20152# vss nfet$247
Xnfet$273_0 m1_n8283_20611# vss m1_n8283_19850# vss nfet$273
Xpfet$258_0 vdd vdd vdd m1_n5019_19550# m1_n4485_20152# m1_n4485_20152# pfet$258
Xnfet$242_82 m1_11415_25662# m1_12259_24224# m1_13363_25658# vss nfet$242
Xnfet$242_71 m1_28147_25662# m1_28371_23922# m1_28635_24542# vss nfet$242
Xnfet$242_60 pd6 vss m1_16322_21786# vss nfet$242
Xnfet$245_4 m1_10299_17343# m1_10560_16202# m1_10075_17518# vss nfet$245
Xnfet$247_16 m1_17381_17714# vss m1_19969_19550# vss nfet$247
Xpfet$251_7 vdd vdd m1_n10452_25858# m1_n4978_24224# pfet$251
Xpfet$235_11 vdd vdd m1_32817_25662# m1_32675_25947# pfet$235
Xpfet$227_100 vdd vdd m1_29607_24346# m1_n7513_20152# pfet$227
Xnfet$243_1 m1_n1263_21786# m1_n1263_21786# m1_354_22513# m1_354_22513# m1_n42_21586#
+ vss nfet$243
Xnfet$250_2 m1_n1271_25858# vss m1_n1134_25662# vss nfet$250
Xpfet$228_1 vdd vdd m1_11381_15778# m1_11738_16080# pfet$228
Xpfet$235_2 vdd vdd m1_n1271_25858# m1_n10452_25858# pfet$235
Xnfet$244_17 m1_12935_19550# m1_12935_19550# vss vss m1_13373_20470# vss nfet$244
Xpfet$240_0 vdd vdd m1_n1263_21786# pd1 pfet$240
Xpfet$232_12 vdd vdd m1_26676_16080# m1_n7513_20152# pfet$232
Xnfet$245_82 m1_10299_17343# vss m1_10458_17836# vss nfet$245
Xnfet$245_71 m1_14641_17836# m1_15921_16080# m1_15454_18030# vss nfet$245
Xnfet$245_60 m1_18665_17343# vss m1_18824_17836# vss nfet$245
Xpfet$227_89 vdd vdd m1_19839_21786# pd7 pfet$227
Xpfet$227_78 vdd m1_20269_24542# vdd m1_21241_24346# pfet$227
Xpfet$227_67 vdd m1_15822_23922# m1_16086_24542# m1_15461_25858# pfet$227
Xpfet$227_56 vdd m1_24808_24224# m1_25912_25658# m1_23827_25858# pfet$227
Xpfet$227_45 vdd vdd m1_16442_24224# m1_15822_23922# pfet$227
Xpfet$227_34 vdd m1_9180_25658# m1_9973_24542# m1_7232_25662# pfet$227
Xpfet$227_23 vdd m1_3537_24542# vdd m1_4509_24346# pfet$227
Xpfet$227_12 vdd m1_7577_25858# vdd m1_9180_25658# pfet$227
Xnfet$268_3 m1_n6973_21481# m1_n6973_21481# m1_n6839_20152# m1_n6839_20152# m1_n6282_20470#
+ vss nfet$268
Xnfet$241_18 m1_21241_24346# m1_21241_24346# vss vss m1_20723_24542# vss nfet$241
Xnfet$254_9 m1_25107_21786# m1_25107_21786# vss vss m1_23945_21586# vss nfet$254
Xnfet$273_1 m1_n7513_20152# m1_n8283_19850# vss vss nfet$273
Xnfet$247_8 m1_n7383_17599# vss m1_n1133_19550# vss nfet$247
Xnfet$266_0 m1_n10452_25858# m1_n10452_25858# m1_n7186_25858# m1_n7186_25858# m1_n6629_25502#
+ vss nfet$266
Xnfet$242_72 m1_23827_25858# m1_25912_25658# m1_26705_24542# vss nfet$242
Xnfet$242_61 m1_23964_25662# m1_24808_24224# m1_25912_25658# vss nfet$242
Xnfet$242_50 m1_n7513_20152# vss m1_21241_24346# vss nfet$242
Xnfet$245_5 m1_10458_17836# m1_11738_16080# m1_11271_18030# vss nfet$245
Xnfet$247_17 m1_21880_15478# vss m1_25722_20152# vss nfet$247
Xpfet$235_12 vdd vdd m1_32193_25858# m1_25107_21786# pfet$235
Xpfet$227_101 vdd vdd m1_28010_25858# m1_21590_21786# pfet$227
Xnfet$243_2 m1_9288_21786# m1_9288_21786# m1_9645_21447# m1_9645_21447# m1_10509_21586#
+ vss nfet$243
Xnfet$250_3 m1_n7513_20152# vss m1_326_24346# vss nfet$250
Xpfet$235_3 vdd vdd m1_1607_24542# m1_n789_25858# pfet$235
Xpfet$228_2 vdd m1_12355_15778# m1_11738_16080# m1_10458_17836# pfet$228
Xpfet$240_1 vdd vdd m1_2254_21786# pd2 pfet$240
Xpfet$233_0 vdd vdd m1_2384_19550# m1_n3534_17714# pfet$233
Xpfet$232_13 vdd vdd m1_25747_17714# m1_26217_17714# pfet$232
Xpfet$227_79 vdd m1_17546_25658# m1_18339_24542# m1_15598_25662# pfet$227
Xpfet$227_68 vdd vdd m1_16086_24542# m1_16442_24224# pfet$227
Xpfet$227_57 vdd vdd m1_24451_25662# m1_24309_25858# pfet$227
Xpfet$227_46 vdd m1_16442_24224# m1_17546_25658# m1_15461_25858# pfet$227
Xnfet$245_72 m1_17851_17714# vss m1_18441_17518# vss nfet$245
Xnfet$245_61 m1_20104_16080# vss m1_19747_15778# vss nfet$245
Xnfet$245_50 m1_25747_17714# vss m1_22848_17343# vss nfet$245
Xpfet$227_35 vdd m1_7720_24542# vdd m1_8692_24346# pfet$227
Xpfet$227_24 vdd vdd m1_5790_24542# m1_3394_25858# pfet$227
Xpfet$227_13 vdd vdd m1_12259_24224# m1_11639_23922# pfet$227
Xnfet$268_4 m1_2590_19404# m1_2590_19404# vss vss m1_n2445_21430# vss nfet$268
Xnfet$241_19 m1_21729_25658# m1_21729_25658# vss vss m1_22188_25502# vss nfet$241
Xnfet$247_9 m1_25747_17714# vss m1_27003_19550# vss nfet$247
Xnfet$259_0 m1_34093_22102# vss fout vss nfet$259
Xnfet$273_2 m1_n8145_21908# vss m1_n8283_20611# vss nfet$273
Xnfet$266_1 m1_n6111_25858# m1_n6111_25858# vss vss m1_n6629_25502# vss nfet$266
Xnfet$242_73 m1_24309_25858# vss m1_21590_21786# vss nfet$242
Xnfet$242_62 m1_24188_23922# vss m1_24808_24224# vss nfet$242
Xnfet$242_51 m1_19644_25858# m1_21729_25658# m1_22522_24542# vss nfet$242
Xnfet$242_40 m1_15598_25662# m1_16442_24224# m1_17546_25658# vss nfet$242
Xnfet$245_6 m1_6116_17343# vss m1_6275_17836# vss nfet$245
Xpfet$235_13 vdd vdd m1_33790_24346# m1_n7513_20152# pfet$235
Xpfet$227_102 vdd m1_28371_23922# m1_28635_24542# m1_28010_25858# pfet$227
Xnfet$243_3 m1_9418_21590# m1_9418_21590# m1_9645_21447# m1_9645_21447# m1_9877_21586#
+ vss nfet$243
Xnfet$250_4 m1_n789_25858# vss m1_1607_24542# vss nfet$250
Xpfet$235_4 vdd vdd m1_488_21786# m1_n789_25858# pfet$235
Xpfet$228_3 vdd m1_11381_15778# m1_10560_16202# m1_10299_17343# pfet$228
Xnfet$241_0 m1_4509_24346# m1_4509_24346# vss vss m1_3991_24542# vss nfet$241
Xpfet$240_2 vdd vdd m1_26873_21786# pd9 pfet$240
Xpfet$233_1 vdd vdd m1_4620_20152# m1_n3218_15478# pfet$233
Xpfet$227_69 vdd vdd m1_12875_24346# m1_n7513_20152# pfet$227
Xpfet$227_58 vdd vdd m1_23964_25662# m1_23827_25858# pfet$227
Xpfet$227_47 vdd vdd m1_15943_25858# m1_17058_24346# pfet$227
Xnfet$245_73 m1_13668_17714# vss m1_16538_15778# vss nfet$245
Xnfet$245_62 m1_18665_17343# m1_20721_15778# m1_20104_16080# vss nfet$245
Xnfet$245_51 m1_n7513_20152# vss m1_22493_16080# vss nfet$245
Xpfet$227_36 vdd vdd m1_8692_24346# m1_n7513_20152# pfet$227
Xpfet$227_25 vdd vdd m1_4005_21786# m1_3394_25858# pfet$227
Xpfet$227_14 vdd vdd m1_11902_25662# m1_11760_25858# pfet$227
Xnfet$245_40 m1_n2250_17343# m1_n194_15778# m1_n811_16080# vss nfet$245
Xnfet$268_5 m1_6107_19404# m1_6107_19404# m1_n5227_21418# m1_n5227_21418# m1_n2445_21430#
+ vss nfet$268
Xnfet$273_3 m1_n8283_19850# m1_n8283_20611# vss vss nfet$273
Xnfet$242_63 m1_14556_21786# vss m1_19644_25858# vss nfet$242
Xnfet$242_52 m1_20126_25858# vss m1_22522_24542# vss nfet$242
Xnfet$242_41 pd5 vss m1_12805_21786# vss nfet$242
Xnfet$242_30 m1_n7513_20152# vss m1_17058_24346# vss nfet$242
Xpfet$228_90 vdd m1_19747_15778# m1_18926_16202# m1_18665_17343# pfet$228
Xnfet$242_74 pd8 vss m1_23356_21786# vss nfet$242
Xnfet$245_7 m1_9485_17714# vss m1_10075_17518# vss nfet$245
Xpfet$256_0 vdd m1_n6380_21786# m1_n6380_21786# m1_n5019_19550# m1_n5227_20152# m1_n5227_20152#
+ pfet$256
Xnfet$271_0 m1_n10933_25858# m1_n8848_25658# m1_n8055_24542# vss nfet$271
Xpfet$227_103 vdd vdd m1_28635_24542# m1_28991_24224# pfet$227
Xnfet$250_5 m1_n789_25858# vss m1_488_21786# vss nfet$250
Xpfet$235_5 vdd vdd m1_326_24346# m1_n7513_20152# pfet$235
Xpfet$228_4 vdd m1_9485_17714# vdd m1_10560_16202# pfet$228
Xnfet$243_4 m1_5901_21590# m1_5901_21590# m1_7388_22513# m1_7388_22513# m1_6360_21586#
+ vss nfet$243
Xnfet$241_1 m1_3893_24224# m1_3893_24224# m1_3537_24542# m1_3537_24542# m1_3991_24542#
+ vss nfet$241
Xpfet$233_2 vdd vdd m1_1103_20152# m1_n7401_15478# pfet$233
Xpfet$227_59 vdd vdd m1_16322_21786# pd6 pfet$227
Xpfet$227_48 vdd m1_16085_25662# m1_15822_23922# m1_15598_25662# pfet$227
Xnfet$245_74 m1_14482_17343# vss m1_14641_17836# vss nfet$245
Xnfet$245_63 m1_13668_17714# vss m1_14258_17518# vss nfet$245
Xnfet$245_52 m1_23007_17836# m1_24287_16080# m1_23820_18030# vss nfet$245
Xpfet$227_37 vdd vdd m1_9973_24542# m1_7577_25858# pfet$227
Xpfet$227_26 vdd m1_4997_25658# m1_5790_24542# m1_3049_25662# pfet$227
Xpfet$227_15 vdd m1_11902_25662# m1_11639_23922# m1_11415_25662# pfet$227
Xnfet$245_30 sd6 vss m1_5148_15478# vss nfet$245
Xnfet$245_41 m1_n2091_17836# m1_n1168_15778# m1_n1989_16202# vss nfet$245
Xnfet$268_6 m1_n5764_21786# m1_n5764_21786# vss vss m1_n6282_21430# vss nfet$268
Xpfet$228_91 vdd m1_24287_16080# m1_23820_18030# m1_22848_17343# pfet$228
Xpfet$228_80 vdd vdd m1_15564_15778# m1_15921_16080# pfet$228
Xnfet$242_75 m1_28371_23922# vss m1_28991_24224# vss nfet$242
Xnfet$242_64 m1_19644_25858# vss m1_19781_25662# vss nfet$242
Xnfet$242_53 m1_23827_25858# m1_24451_25662# m1_24188_23922# vss nfet$242
Xnfet$242_42 m1_15943_25858# vss m1_16085_25662# vss nfet$242
Xnfet$242_31 m1_15943_25858# vss m1_18339_24542# vss nfet$242
Xnfet$242_20 pd3 vss m1_5771_21786# vss nfet$242
Xnfet$245_8 m1_7555_16080# vss m1_7198_15778# vss nfet$245
Xnfet$264_0 m1_n6274_17836# m1_n4994_16080# m1_n5461_18030# vss nfet$264
Xnfet$271_1 m1_n10796_25662# m1_n10572_23922# m1_n10308_24542# vss nfet$271
Xpfet$256_1 vdd vdd vdd m1_n5019_22344# m1_n4485_21904# m1_n4485_21904# pfet$256
Xpfet$249_0 vdd m1_n10309_25662# m1_n10572_23922# m1_n10796_25662# pfet$249
Xpfet$227_104 vdd m1_25912_25658# m1_26705_24542# m1_23964_25662# pfet$227
Xnfet$250_6 m1_n910_23922# vss m1_n290_24224# vss nfet$250
Xpfet$235_6 vdd vdd m1_n290_24224# m1_n910_23922# pfet$235
Xnfet$243_5 m1_2254_21786# m1_2254_21786# m1_3871_22513# m1_3871_22513# m1_3475_21586#
+ vss nfet$243
Xpfet$228_5 vdd m1_7198_15778# m1_6377_16202# m1_6116_17343# pfet$228
Xnfet$241_2 m1_4997_25658# m1_4997_25658# vss vss m1_5456_25502# vss nfet$241
Xpfet$233_3 vdd vdd m1_5901_19550# m1_649_17714# pfet$233
Xnfet$245_75 sd3 vss m1_17697_15478# vss nfet$245
Xnfet$245_64 m1_13668_17714# vss m1_13198_17714# vss nfet$245
Xnfet$245_53 m1_22848_17343# vss m1_23007_17836# vss nfet$245
Xnfet$245_31 m1_1933_17343# m1_3989_15778# m1_3372_16080# vss nfet$245
Xnfet$245_20 m1_1119_17714# vss m1_1709_17518# vss nfet$245
Xnfet$245_42 m1_n811_16080# vss m1_n1168_15778# vss nfet$245
Xpfet$231_0 vdd vdd m1_n1133_21590# m1_n1263_21786# pfet$231
Xpfet$227_49 vdd m1_20126_25858# vdd m1_21729_25658# pfet$227
Xpfet$227_38 vdd vdd m1_16085_25662# m1_15943_25858# pfet$227
Xpfet$227_27 vdd vdd m1_11278_25858# m1_7522_21786# pfet$227
Xpfet$227_16 vdd vdd m1_5771_21786# pd3 pfet$227
Xnfet$268_7 m1_n3822_21786# m1_n3822_21786# m1_n4485_21904# m1_n4485_21904# m1_n3724_21430#
+ vss nfet$268
Xpfet$228_92 vdd m1_15454_18030# vdd m1_14127_16080# pfet$228
Xpfet$228_81 vdd vdd m1_13668_17714# m1_14127_16080# pfet$228
Xpfet$228_70 vdd vdd m1_18824_17836# m1_18665_17343# pfet$228
Xnfet$242_76 m1_28492_25858# vss m1_28634_25662# vss nfet$242
Xnfet$242_65 m1_28492_25858# vss m1_25107_21786# vss nfet$242
Xnfet$242_54 m1_24309_25858# vss m1_24451_25662# vss nfet$242
Xnfet$242_43 m1_15461_25858# vss m1_15598_25662# vss nfet$242
Xnfet$242_32 m1_15461_25858# m1_17546_25658# m1_18339_24542# vss nfet$242
Xnfet$242_21 m1_11278_25858# m1_11902_25662# m1_11639_23922# vss nfet$242
Xnfet$242_10 m1_7577_25858# vss m1_9973_24542# vss nfet$242
Xnfet$245_9 sd5 vss m1_9331_15478# vss nfet$245
Xnfet$257_0 m1_31535_22102# m1_32818_21586# vss vss nfet$257
Xnfet$264_1 m1_n6433_17343# m1_n4377_15778# m1_n4994_16080# vss nfet$264
Xnfet$271_2 m1_n10933_25858# m1_n10309_25662# m1_n10572_23922# vss nfet$271
Xpfet$256_2 vdd m1_n5764_21786# m1_n5764_21786# m1_n5019_22344# m1_n5227_21418# m1_n5227_21418#
+ pfet$256
Xpfet$249_1 vdd m1_n9952_24224# m1_n8848_25658# m1_n10933_25858# pfet$249
Xpfet$227_105 vdd vdd m1_30888_24542# m1_28492_25858# pfet$227
Xnfet$250_7 m1_25107_21786# vss m1_32193_25858# vss nfet$250
Xnfet$243_6 m1_2384_21590# m1_2384_21590# m1_3871_22513# m1_3871_22513# m1_2843_21586#
+ vss nfet$243
Xpfet$235_7 vdd vdd m1_32330_25662# m1_32193_25858# pfet$235
Xpfet$228_6 vdd vdd m1_7198_15778# m1_7555_16080# pfet$228
Xnfet$241_3 m1_4509_24346# m1_4509_24346# m1_3394_25858# m1_3394_25858# m1_5456_25502#
+ vss nfet$241
Xpfet$233_4 vdd vdd m1_12935_19550# m1_9015_17714# pfet$233
Xnfet$250_10 m1_32675_25947# vss m1_35071_24542# vss nfet$250
Xnfet$245_76 m1_14482_17343# m1_16538_15778# m1_15921_16080# vss nfet$245
Xnfet$245_65 m1_14482_17343# m1_14743_16202# m1_14258_17518# vss nfet$245
Xnfet$245_54 m1_22848_17343# m1_23109_16202# m1_22624_17518# vss nfet$245
Xnfet$245_32 m1_2092_17836# m1_3015_15778# m1_2194_16202# vss nfet$245
Xnfet$245_21 m1_1933_17343# m1_2194_16202# m1_1709_17518# vss nfet$245
Xnfet$245_10 m1_11738_16080# vss m1_11381_15778# vss nfet$245
Xnfet$245_43 sd8 vss m1_n3218_15478# vss nfet$245
Xpfet$231_1 vdd vdd m1_11671_21786# m1_11039_21786# pfet$231
Xpfet$227_39 vdd vdd m1_15598_25662# m1_15461_25858# pfet$227
Xnfet$261_20 m1_22493_16080# m1_22493_16080# m1_22034_17714# m1_22034_17714# m1_22591_16398#
+ vss nfet$261
Xpfet$227_28 vdd m1_11639_23922# m1_11903_24542# m1_11278_25858# pfet$227
Xpfet$227_17 vdd vdd m1_7577_25858# m1_8692_24346# pfet$227
Xnfet$268_8 m1_9624_19404# m1_9624_19404# vss vss m1_n3724_21430# vss nfet$268
Xpfet$228_93 vdd m1_23820_18030# vdd m1_22493_16080# pfet$228
Xpfet$228_82 vdd m1_13668_17714# vdd m1_14743_16202# pfet$228
Xpfet$228_71 vdd vdd m1_19747_15778# m1_20104_16080# pfet$228
Xpfet$228_60 vdd vdd m1_n194_15778# m1_n3064_17714# pfet$228
Xnfet$242_77 m1_28010_25858# vss m1_28147_25662# vss nfet$242
Xnfet$242_66 m1_28010_25858# m1_30095_25658# m1_30888_24542# vss nfet$242
Xnfet$242_55 m1_23827_25858# vss m1_23964_25662# vss nfet$242
Xnfet$242_44 m1_15822_23922# vss m1_16442_24224# vss nfet$242
Xnfet$242_33 m1_11760_25858# vss m1_14156_24542# vss nfet$242
Xnfet$242_22 m1_11760_25858# vss m1_11902_25662# vss nfet$242
Xnfet$242_11 m1_7522_21786# vss m1_11278_25858# vss nfet$242
Xnfet$264_2 m1_n6274_17836# m1_n5351_15778# m1_n6172_16202# vss nfet$264
Xnfet$271_3 m1_n10796_25662# m1_n9952_24224# m1_n8848_25658# vss nfet$271
Xpfet$249_2 vdd m1_n4362_24346# m1_n4847_25662# m1_n4464_25980# pfet$249
Xpfet$227_106 vdd vdd m1_25107_21786# m1_28492_25858# pfet$227
Xnfet$250_8 m1_32193_25858# vss m1_32330_25662# vss nfet$250
Xnfet$243_7 m1_5771_21786# m1_5771_21786# m1_7388_22513# m1_7388_22513# m1_6992_21586#
+ vss nfet$243
Xpfet$235_8 vdd vdd m1_33174_24224# m1_32554_23922# pfet$235
Xpfet$228_7 vdd vdd m1_6275_17836# m1_6116_17343# pfet$228
Xpfet$254_0 vdd vdd m1_n7186_25858# m1_n10452_25858# pfet$254
Xnfet$241_4 m1_12259_24224# m1_12259_24224# m1_11903_24542# m1_11903_24542# m1_12357_24542#
+ vss nfet$241
Xpfet$233_5 vdd vdd m1_8137_20152# m1_965_15478# pfet$233
Xnfet$250_11 m1_32554_23922# vss m1_33174_24224# vss nfet$250
Xpfet$231_2 vdd vdd m1_12935_21590# m1_12805_21786# pfet$231
Xnfet$245_77 sd4 vss m1_13514_15478# vss nfet$245
Xnfet$245_66 m1_n7513_20152# vss m1_14127_16080# vss nfet$245
Xnfet$261_21 m1_14127_16080# m1_14127_16080# vss vss m1_15690_17358# vss nfet$261
Xnfet$245_55 m1_22034_17714# vss m1_24904_15778# vss nfet$245
Xnfet$245_44 m1_n2091_17836# m1_n811_16080# m1_n1278_18030# vss nfet$245
Xpfet$227_29 vdd vdd m1_11903_24542# m1_12259_24224# pfet$227
Xpfet$227_18 vdd vdd m1_11415_25662# m1_11278_25858# pfet$227
Xnfet$245_33 sd7 vss m1_965_15478# vss nfet$245
Xnfet$261_10 m1_1578_16080# m1_1578_16080# m1_1119_17714# m1_1119_17714# m1_1676_16398#
+ vss nfet$261
Xnfet$245_22 m1_6116_17343# m1_6377_16202# m1_5892_17518# vss nfet$245
Xnfet$245_11 m1_10299_17343# m1_12355_15778# m1_11738_16080# vss nfet$245
Xnfet$268_9 m1_n6380_21786# m1_n6380_21786# m1_n6839_21786# m1_n6839_21786# m1_n6282_21430#
+ vss nfet$268
Xnfet$242_78 m1_28010_25858# m1_28634_25662# m1_28371_23922# vss nfet$242
Xnfet$242_67 m1_28492_25858# vss m1_30888_24542# vss nfet$242
Xnfet$242_56 m1_19781_25662# m1_20625_24224# m1_21729_25658# vss nfet$242
Xnfet$242_45 m1_15461_25858# m1_16085_25662# m1_15822_23922# vss nfet$242
Xnfet$242_34 m1_11278_25858# m1_13363_25658# m1_14156_24542# vss nfet$242
Xpfet$228_94 vdd vdd m1_22624_17518# m1_22034_17714# pfet$228
Xpfet$228_83 vdd m1_16538_15778# m1_15921_16080# m1_14641_17836# pfet$228
Xpfet$228_72 vdd m1_20721_15778# m1_20104_16080# m1_18824_17836# pfet$228
Xpfet$228_61 vdd m1_n811_16080# m1_n1278_18030# m1_n2250_17343# pfet$228
Xnfet$242_23 m1_11278_25858# vss m1_11415_25662# vss nfet$242
Xnfet$242_12 m1_7577_25858# vss m1_7522_21786# vss nfet$242
Xpfet$228_50 vdd m1_n1168_15778# m1_n1989_16202# m1_n2250_17343# pfet$228
Xnfet$264_3 m1_n6433_17343# m1_n6172_16202# m1_n6657_17518# vss nfet$264
Xnfet$271_4 m1_n4623_25487# m1_n2567_23922# m1_n3184_24224# vss nfet$271
Xpfet$249_3 vdd m1_n3184_24224# m1_n3651_26174# m1_n4623_25487# pfet$249
Xpfet$227_107 vdd m1_24309_25858# vdd m1_25912_25658# pfet$227
Xnfet$250_9 m1_n7513_20152# vss m1_33790_24346# vss nfet$250
Xnfet$243_8 m1_23486_21590# m1_23486_21590# m1_24973_22513# m1_24973_22513# m1_23945_21586#
+ vss nfet$243
Xpfet$235_9 vdd vdd m1_28624_21786# m1_32675_25947# pfet$235
Xnfet$262_0 m1_4620_20152# m1_4620_20152# m1_2590_19404# m1_2590_19404# m1_3454_20470#
+ vss nfet$262
Xpfet$228_8 vdd vdd m1_9331_15478# sd5 pfet$228
Xpfet$247_0 vdd vdd m1_n7513_20152# m1_35837_22102# pfet$247
Xpfet$254_1 vdd m1_n7186_25858# vdd m1_n6111_25858# pfet$254
Xnfet$241_5 m1_8692_24346# m1_8692_24346# vss vss m1_8174_24542# vss nfet$241
Xnfet$250_12 m1_32675_25947# vss m1_28624_21786# vss nfet$250
Xpfet$233_6 vdd vdd m1_9418_19550# m1_4832_17714# pfet$233
Xpfet$231_3 vdd vdd m1_9418_21590# m1_9288_21786# pfet$231
Xnfet$245_78 m1_14641_17836# m1_15564_15778# m1_14743_16202# vss nfet$245
Xnfet$261_22 m1_15564_15778# m1_15564_15778# m1_15454_18030# m1_15454_18030# m1_15690_17358#
+ vss nfet$261
Xnfet$245_67 m1_17381_17714# vss m1_14482_17343# vss nfet$245
Xnfet$245_56 m1_24287_16080# vss m1_23930_15778# vss nfet$245
Xnfet$245_45 m1_n3064_17714# vss m1_n194_15778# vss nfet$245
Xpfet$227_19 vdd vdd m1_7095_25858# m1_4005_21786# pfet$227
Xnfet$245_34 m1_n2250_17343# vss m1_n2091_17836# vss nfet$245
Xnfet$245_23 m1_5302_17714# vss m1_4832_17714# vss nfet$245
Xnfet$245_12 m1_9485_17714# vss m1_12355_15778# vss nfet$245
Xnfet$261_11 m1_6377_16202# m1_6377_16202# vss vss m1_5859_16398# vss nfet$261
Xnfet$242_79 pd7 vss m1_19839_21786# vss nfet$242
Xnfet$242_68 m1_n7513_20152# vss m1_29607_24346# vss nfet$242
Xnfet$242_57 m1_20126_25858# vss m1_20268_25662# vss nfet$242
Xnfet$242_46 m1_20126_25858# vss m1_18073_21786# vss nfet$242
Xnfet$242_35 m1_15598_25662# m1_15822_23922# m1_16086_24542# vss nfet$242
Xpfet$228_95 vdd vdd m1_21564_17714# m1_22034_17714# pfet$228
Xpfet$228_84 vdd vdd m1_17381_17714# m1_17851_17714# pfet$228
Xpfet$228_73 vdd vdd m1_16538_15778# m1_13668_17714# pfet$228
Xpfet$228_62 vdd vdd m1_23007_17836# m1_22848_17343# pfet$228
Xnfet$242_24 m1_7095_25858# m1_7719_25662# m1_7456_23922# vss nfet$242
Xnfet$242_13 m1_11415_25662# m1_11639_23922# m1_11903_24542# vss nfet$242
Xpfet$228_40 vdd m1_10560_16202# m1_10075_17518# m1_10458_17836# pfet$228
Xpfet$228_51 vdd vdd m1_n1168_15778# m1_n811_16080# pfet$228
Xpfet$230_30 vdd vdd vdd m1_24560_19550# m1_21880_15478# m1_21880_15478# pfet$230
Xnfet$264_4 m1_27031_17343# m1_27292_16202# m1_26807_17518# vss nfet$264
Xnfet$271_5 m1_n4464_25980# m1_n3541_23922# m1_n4362_24346# vss nfet$271
Xpfet$249_4 vdd m1_n2567_23922# m1_n3184_24224# m1_n4464_25980# pfet$249
Xpfet$227_108 vdd vdd m1_25424_24346# m1_n7513_20152# pfet$227
Xnfet$243_9 m1_23356_21786# m1_23356_21786# m1_24973_22513# m1_24973_22513# m1_24577_21586#
+ vss nfet$243
Xnfet$255_0 m1_21456_22513# m1_21456_22513# m1_30256_19792# m1_30256_19792# m1_30492_20470#
+ vss nfet$255
Xnfet$262_1 m1_1103_20152# m1_1103_20152# m1_n927_19404# m1_n927_19404# m1_n63_20470#
+ vss nfet$262
Xpfet$228_9 vdd vdd m1_8172_15778# m1_5302_17714# pfet$228
Xnfet$241_6 m1_8076_24224# m1_8076_24224# m1_7720_24542# m1_7720_24542# m1_8174_24542#
+ vss nfet$241
Xpfet$233_7 vdd vdd m1_11654_20152# m1_5148_15478# pfet$233
Xnfet$250_13 m1_32675_25947# vss m1_32817_25662# vss nfet$250
Xnfet$245_79 m1_15921_16080# vss m1_15564_15778# vss nfet$245
Xnfet$261_23 m1_18926_16202# m1_18926_16202# vss vss m1_18408_16398# vss nfet$261
Xnfet$245_68 m1_18665_17343# m1_18926_16202# m1_18441_17518# vss nfet$245
Xnfet$245_57 m1_22848_17343# m1_24904_15778# m1_24287_16080# vss nfet$245
Xnfet$245_46 m1_22034_17714# vss m1_21564_17714# vss nfet$245
Xnfet$245_24 m1_4832_17714# vss m1_1933_17343# vss nfet$245
Xnfet$245_13 m1_10458_17836# m1_11381_15778# m1_10560_16202# vss nfet$245
Xnfet$245_35 m1_n7513_20152# vss m1_5761_16080# vss nfet$245
Xnfet$261_12 m1_n1168_15778# m1_n1168_15778# m1_n1278_18030# m1_n1278_18030# m1_n1042_17358#
+ vss nfet$261
Xpfet$231_4 vdd vdd m1_8154_21786# m1_7522_21786# pfet$231
Xpfet$228_96 vdd vdd m1_18665_17343# m1_21564_17714# pfet$228
Xpfet$228_85 vdd m1_18926_16202# m1_18441_17518# m1_18824_17836# pfet$228
Xpfet$228_74 vdd vdd m1_14641_17836# m1_14482_17343# pfet$228
Xpfet$228_63 vdd m1_23930_15778# m1_23109_16202# m1_22848_17343# pfet$228
Xpfet$228_30 vdd vdd m1_1933_17343# m1_4832_17714# pfet$228
Xpfet$228_41 vdd vdd m1_10075_17518# m1_9485_17714# pfet$228
Xpfet$228_52 vdd m1_n3064_17714# vdd m1_n1989_16202# pfet$228
Xnfet$242_69 m1_24309_25858# vss m1_26705_24542# vss nfet$242
Xnfet$242_58 m1_20005_23922# vss m1_20625_24224# vss nfet$242
Xnfet$242_47 m1_23964_25662# m1_24188_23922# m1_24452_24542# vss nfet$242
Xnfet$242_36 m1_11760_25858# vss m1_11039_21786# vss nfet$242
Xnfet$242_25 m1_7232_25662# m1_8076_24224# m1_9180_25658# vss nfet$242
Xnfet$242_14 m1_n7513_20152# vss m1_8692_24346# vss nfet$242
Xpfet$230_31 vdd m1_n2543_20130# m1_n2543_20130# m1_20407_19850# m1_19969_19550# m1_19969_19550#
+ pfet$230
Xpfet$230_20 vdd m1_n3822_21786# m1_n3822_21786# m1_14009_19550# m1_9015_17714# m1_9015_17714#
+ pfet$230
Xnfet$264_5 m1_27031_17343# m1_29087_15778# m1_28470_16080# vss nfet$264
Xnfet$271_6 m1_n4464_25980# m1_n3184_24224# m1_n3651_26174# vss nfet$271
Xpfet$249_5 vdd m1_n10572_23922# m1_n10308_24542# m1_n10933_25858# pfet$249
Xpfet$227_109 vdd m1_12259_24224# m1_13363_25658# m1_11278_25858# pfet$227
Xnfet$262_2 m1_n3218_15478# m1_n3218_15478# m1_2590_19404# m1_2590_19404# m1_2822_20470#
+ vss nfet$262
Xnfet$255_1 m1_14422_22513# m1_14422_22513# m1_31535_19792# m1_31535_19792# m1_31771_20470#
+ vss nfet$255
Xnfet$248_0 sd9 vss m1_n7401_15478# vss nfet$248
Xnfet$241_7 m1_9180_25658# m1_9180_25658# vss vss m1_9639_25502# vss nfet$241
Xpfet$233_8 vdd vdd m1_n1133_19550# m1_n7383_17599# pfet$233
Xpfet$252_0 vdd vdd m1_n4485_20152# m1_n3822_20130# pfet$252
Xnfet$261_24 m1_18310_16080# m1_18310_16080# m1_17851_17714# m1_17851_17714# m1_18408_16398#
+ vss nfet$261
Xnfet$245_69 m1_17851_17714# vss m1_17381_17714# vss nfet$245
Xnfet$245_58 m1_23007_17836# m1_23930_15778# m1_23109_16202# vss nfet$245
Xnfet$245_47 m1_22034_17714# vss m1_22624_17518# vss nfet$245
Xnfet$245_25 m1_2092_17836# m1_3372_16080# m1_2905_18030# vss nfet$245
Xnfet$245_14 m1_6116_17343# m1_8172_15778# m1_7555_16080# vss nfet$245
Xnfet$245_36 m1_n3064_17714# vss m1_n2474_17518# vss nfet$245
Xnfet$261_13 m1_n2605_16080# m1_n2605_16080# vss vss m1_n1042_17358# vss nfet$261
Xpfet$231_5 vdd vdd m1_1120_21786# m1_488_21786# pfet$231
Xpfet$228_97 vdd vdd m1_22493_16080# m1_n7513_20152# pfet$228
Xpfet$228_86 vdd m1_19637_18030# vdd m1_18310_16080# pfet$228
Xpfet$228_75 vdd vdd m1_17697_15478# sd3 pfet$228
Xpfet$228_64 vdd vdd m1_23930_15778# m1_24287_16080# pfet$228
Xpfet$228_20 vdd vdd m1_1119_17714# m1_1578_16080# pfet$228
Xpfet$228_31 vdd m1_3372_16080# m1_2905_18030# m1_1933_17343# pfet$228
Xpfet$228_42 vdd m1_11271_18030# vdd m1_9944_16080# pfet$228
Xpfet$228_53 vdd vdd m1_n3218_15478# sd8 pfet$228
Xnfet$242_59 m1_19644_25858# m1_20268_25662# m1_20005_23922# vss nfet$242
Xnfet$242_48 m1_18073_21786# vss m1_23827_25858# vss nfet$242
Xnfet$242_37 m1_11039_21786# vss m1_15461_25858# vss nfet$242
Xnfet$242_26 m1_7095_25858# m1_9180_25658# m1_9973_24542# vss nfet$242
Xnfet$242_15 m1_7232_25662# m1_7456_23922# m1_7720_24542# vss nfet$242
Xpfet$230_32 vdd m1_n2543_20130# m1_n2543_20130# m1_21043_19550# m1_17381_17714# m1_17381_17714#
+ pfet$230
Xpfet$230_21 vdd vdd vdd m1_13373_19850# m1_15171_20152# m1_15171_20152# pfet$230
Xnfet$264_6 m1_27190_17836# m1_28113_15778# m1_27292_16202# vss nfet$264
Xpfet$230_10 vdd vdd vdd m1_9856_19850# m1_11654_20152# m1_11654_20152# pfet$230
Xnfet$271_7 m1_n4623_25487# m1_n4362_24346# m1_n4847_25662# vss nfet$271
Xpfet$249_6 vdd m1_n8848_25658# m1_n8055_24542# m1_n10796_25662# pfet$249
Xnfet$248_1 sd2 vss m1_21880_15478# vss nfet$248
Xnfet$255_2 m1_17939_22513# m1_17939_22513# vss vss m1_31771_20470# vss nfet$255
Xnfet$262_3 m1_8137_20152# m1_8137_20152# m1_6107_19404# m1_6107_19404# m1_6971_20470#
+ vss nfet$262
Xnfet$260_0 fout vss m1_35837_22102# vss nfet$260
Xpfet$233_9 vdd vdd m1_27003_19550# m1_25747_17714# pfet$233
Xnfet$241_8 m1_8692_24346# m1_8692_24346# m1_7577_25858# m1_7577_25858# m1_9639_25502#
+ vss nfet$241
Xpfet$245_0 vdd vdd m1_n7247_17714# m1_n6788_16080# pfet$245
Xpfet$252_1 vdd m1_n4485_21904# vdd m1_9624_19404# pfet$252
Xnfet$245_59 m1_17851_17714# vss m1_20721_15778# vss nfet$245
Xnfet$245_48 m1_18824_17836# m1_20104_16080# m1_19637_18030# vss nfet$245
Xnfet$245_26 m1_5302_17714# vss m1_5892_17518# vss nfet$245
Xnfet$245_15 m1_5302_17714# vss m1_8172_15778# vss nfet$245
Xnfet$245_37 m1_n7513_20152# vss m1_n2605_16080# vss nfet$245
Xpfet$231_6 vdd vdd m1_5901_21590# m1_5771_21786# pfet$231
Xnfet$261_25 m1_14743_16202# m1_14743_16202# vss vss m1_14225_16398# vss nfet$261
Xnfet$261_14 m1_n2605_16080# m1_n2605_16080# m1_n3064_17714# m1_n3064_17714# m1_n2507_16398#
+ vss nfet$261
Xpfet$233_10 vdd vdd m1_29239_20152# m1_26063_15478# pfet$233
Xpfet$228_98 vdd m1_20104_16080# m1_19637_18030# m1_18665_17343# pfet$228
Xpfet$228_87 vdd vdd m1_18310_16080# m1_n7513_20152# pfet$228
Xpfet$228_76 vdd m1_17851_17714# vdd m1_18926_16202# pfet$228
Xpfet$228_65 vdd m1_24904_15778# m1_24287_16080# m1_23007_17836# pfet$228
Xpfet$228_21 vdd vdd m1_965_15478# sd7 pfet$228
Xpfet$228_10 vdd m1_8172_15778# m1_7555_16080# m1_6275_17836# pfet$228
Xpfet$228_32 vdd vdd m1_2905_18030# m1_3015_15778# pfet$228
Xpfet$228_43 vdd vdd m1_11271_18030# m1_11381_15778# pfet$228
Xpfet$228_54 vdd vdd m1_n1278_18030# m1_n1168_15778# pfet$228
Xnfet$242_49 m1_19781_25662# m1_20005_23922# m1_20269_24542# vss nfet$242
Xnfet$242_38 m1_n7513_20152# vss m1_12875_24346# vss nfet$242
Xnfet$242_27 m1_7577_25858# vss m1_7719_25662# vss nfet$242
Xnfet$242_16 m1_4005_21786# vss m1_7095_25858# vss nfet$242
Xnfet$264_7 m1_27190_17836# m1_28470_16080# m1_28003_18030# vss nfet$264
Xpfet$230_33 vdd m1_n3206_20274# m1_n3206_20274# m1_24560_19550# m1_21564_17714# m1_21564_17714#
+ pfet$230
Xpfet$230_22 vdd vdd vdd m1_14009_19550# m1_9331_15478# m1_9331_15478# pfet$230
Xpfet$230_11 vdd vdd vdd m1_10492_19550# m1_5148_15478# m1_5148_15478# pfet$230
Xpfet$249_7 vdd m1_n3541_23922# m1_n4362_24346# m1_n4623_25487# pfet$249
Xnfet$248_2 sd1 vss m1_26063_15478# vss nfet$248
Xnfet$255_3 m1_24973_22513# m1_24973_22513# vss vss m1_30492_20470# vss nfet$255
Xnfet$262_4 m1_965_15478# m1_965_15478# m1_6107_19404# m1_6107_19404# m1_6339_20470#
+ vss nfet$262
Xnfet$241_9 m1_17058_24346# m1_17058_24346# vss vss m1_16540_24542# vss nfet$241
Xnfet$260_1 define m1_35837_22102# vss vss nfet$260
Xpfet$238_0 vdd m1_31535_19792# vdd m1_17939_22513# pfet$238
Xpfet$245_1 vdd m1_n7247_17714# vdd m1_n6172_16202# pfet$245
Xpfet$252_2 vdd m1_n5227_21418# vdd m1_2590_19404# pfet$252
Xnfet$253_0 m1_n290_24224# m1_n290_24224# m1_n646_24542# m1_n646_24542# m1_n192_24542#
+ vss nfet$253
Xpfet$231_7 vdd vdd m1_4637_21786# m1_4005_21786# pfet$231
Xnfet$261_26 m1_14127_16080# m1_14127_16080# m1_13668_17714# m1_13668_17714# m1_14225_16398#
+ vss nfet$261
Xnfet$245_49 m1_21564_17714# vss m1_18665_17343# vss nfet$245
Xnfet$245_27 m1_1119_17714# vss m1_3989_15778# vss nfet$245
Xnfet$245_16 m1_6275_17836# m1_7198_15778# m1_6377_16202# vss nfet$245
Xnfet$245_38 m1_n2250_17343# m1_n1989_16202# m1_n2474_17518# vss nfet$245
Xnfet$261_15 m1_n1989_16202# m1_n1989_16202# vss vss m1_n2507_16398# vss nfet$261
Xpfet$233_11 vdd vdd m1_18688_20152# m1_13514_15478# pfet$233
Xpfet$228_22 vdd vdd m1_3015_15778# m1_3372_16080# pfet$228
Xpfet$228_11 vdd vdd m1_9485_17714# m1_9944_16080# pfet$228
Xpfet$228_33 vdd vdd m1_5892_17518# m1_5302_17714# pfet$228
Xnfet$242_39 pd4 vss m1_9288_21786# vss nfet$242
Xpfet$228_99 vdd m1_23109_16202# m1_22624_17518# m1_23007_17836# pfet$228
Xpfet$228_88 vdd vdd m1_18441_17518# m1_17851_17714# pfet$228
Xpfet$228_77 vdd vdd m1_17851_17714# m1_18310_16080# pfet$228
Xpfet$228_66 vdd vdd m1_24904_15778# m1_22034_17714# pfet$228
Xnfet$242_28 m1_3394_25858# vss m1_4005_21786# vss nfet$242
Xnfet$242_17 m1_11639_23922# vss m1_12259_24224# vss nfet$242
Xpfet$228_44 vdd vdd m1_649_17714# m1_1119_17714# pfet$228
Xpfet$228_55 vdd vdd m1_n2474_17518# m1_n3064_17714# pfet$228
Xpfet$230_34 vdd m1_n3206_20274# m1_n3206_20274# m1_23924_19850# m1_23486_19550# m1_23486_19550#
+ pfet$230
Xpfet$230_23 vdd vdd vdd m1_16890_19850# m1_18688_20152# m1_18688_20152# pfet$230
Xpfet$230_12 vdd m1_6107_19404# m1_6107_19404# m1_6975_19550# m1_649_17714# m1_649_17714#
+ pfet$230
Xnfet$255_4 m1_32818_20470# m1_32818_20470# vss vss m1_34329_20470# vss nfet$255
Xnfet$262_5 m1_5148_15478# m1_5148_15478# m1_9624_19404# m1_9624_19404# m1_9856_20470#
+ vss nfet$262
Xnfet$253_1 m1_814_25658# m1_814_25658# vss vss m1_1273_25502# vss nfet$253
Xpfet$245_2 vdd vdd m1_n5461_18030# m1_n5351_15778# pfet$245
Xnfet$246_0 m1_n1263_21786# vss m1_n1133_21590# vss nfet$246
Xpfet$252_3 vdd vdd m1_n5227_21418# m1_6107_19404# pfet$252
Xpfet$238_1 vdd vdd m1_30256_19792# m1_21456_22513# pfet$238
Xpfet$231_8 vdd vdd m1_2384_21590# m1_2254_21786# pfet$231
Xnfet$261_27 m1_18310_16080# m1_18310_16080# vss vss m1_19873_17358# vss nfet$261
Xnfet$261_16 m1_19747_15778# m1_19747_15778# m1_19637_18030# m1_19637_18030# m1_19873_17358#
+ vss nfet$261
Xnfet$245_28 m1_1933_17343# vss m1_2092_17836# vss nfet$245
Xnfet$245_17 m1_649_17714# vss m1_n2250_17343# vss nfet$245
Xnfet$245_39 m1_n3064_17714# vss m1_n3534_17714# vss nfet$245
Xpfet$250_0 vdd vdd m1_n7320_25516# m1_n7186_25858# pfet$250
Xpfet$233_12 vdd vdd m1_15171_20152# m1_9331_15478# pfet$233
Xnfet$242_29 m1_15943_25858# vss m1_14556_21786# vss nfet$242
Xpfet$228_89 vdd vdd m1_22848_17343# m1_25747_17714# pfet$228
Xpfet$228_78 vdd vdd m1_13514_15478# sd4 pfet$228
Xpfet$228_67 vdd m1_22034_17714# vdd m1_23109_16202# pfet$228
Xnfet$242_18 m1_7095_25858# vss m1_7232_25662# vss nfet$242
Xpfet$228_12 vdd m1_3989_15778# m1_3372_16080# m1_2092_17836# pfet$228
Xpfet$228_23 vdd m1_5302_17714# vdd m1_6377_16202# pfet$228
Xpfet$228_34 vdd vdd m1_5761_16080# m1_n7513_20152# pfet$228
Xpfet$228_45 vdd vdd m1_9944_16080# m1_n7513_20152# pfet$228
Xpfet$228_56 vdd m1_n1278_18030# vdd m1_n2605_16080# pfet$228
Xpfet$230_35 vdd m1_n3822_21786# m1_n3822_21786# m1_13373_19850# m1_12935_19550# m1_12935_19550#
+ pfet$230
Xpfet$230_24 vdd m1_n1927_20274# m1_n1927_20274# m1_16890_19850# m1_16452_19550# m1_16452_19550#
+ pfet$230
Xnfet$276_0 m1_n4485_20152# m1_n6380_21786# vss vss nfet$276
Xpfet$230_13 vdd m1_n927_19404# m1_n927_19404# m1_n695_19850# m1_n1133_19550# m1_n1133_19550#
+ pfet$230
Xnfet$255_5 m1_32818_21586# m1_32818_21586# m1_34093_19792# m1_34093_19792# m1_34329_20470#
+ vss nfet$255
Xnfet$262_6 m1_11654_20152# m1_11654_20152# m1_9624_19404# m1_9624_19404# m1_10488_20470#
+ vss nfet$262
Xnfet$253_2 m1_326_24346# m1_326_24346# m1_n789_25858# m1_n789_25858# m1_1273_25502#
+ vss nfet$253
Xnfet$246_1 m1_11039_21786# vss m1_11671_21786# vss nfet$246
Xpfet$238_2 vdd m1_30256_19792# vdd m1_24973_22513# pfet$238
Xpfet$245_3 vdd m1_n5461_18030# vdd m1_n6788_16080# pfet$245
Xpfet$252_4 vdd vdd m1_n4485_21904# m1_n3822_21786# pfet$252
Xpfet$243_0 vdd vdd fout m1_34093_22102# pfet$243
Xpfet$231_9 vdd vdd m1_22222_21786# m1_21590_21786# pfet$231
Xnfet$261_17 m1_22493_16080# m1_22493_16080# vss vss m1_24056_17358# vss nfet$261
Xnfet$245_29 m1_3372_16080# vss m1_3015_15778# vss nfet$245
Xnfet$245_18 m1_1119_17714# vss m1_649_17714# vss nfet$245
Xpfet$250_1 vdd vdd m1_n6111_25858# m1_n6856_24542# pfet$250
Xpfet$233_13 vdd vdd m1_16452_19550# m1_13198_17714# pfet$233
Xpfet$228_79 vdd m1_15564_15778# m1_14743_16202# m1_14482_17343# pfet$228
Xpfet$228_68 vdd vdd m1_22034_17714# m1_22493_16080# pfet$228
Xpfet$228_13 vdd vdd m1_5148_15478# sd6 pfet$228
Xpfet$228_24 vdd m1_6377_16202# m1_5892_17518# m1_6275_17836# pfet$228
Xpfet$228_35 vdd vdd m1_9015_17714# m1_9485_17714# pfet$228
Xpfet$228_46 vdd vdd m1_n2250_17343# m1_649_17714# pfet$228
Xpfet$228_57 vdd m1_n1989_16202# m1_n2474_17518# m1_n2091_17836# pfet$228
Xnfet$242_19 m1_7456_23922# vss m1_8076_24224# vss nfet$242
Xpfet$230_25 vdd vdd vdd m1_17526_19550# m1_13514_15478# m1_13514_15478# pfet$230
Xpfet$230_14 vdd m1_n927_19404# m1_n927_19404# m1_n59_19550# m1_n7383_17599# m1_n7383_17599#
+ pfet$230
Xnfet$276_1 m1_n5227_20152# vss m1_n6380_21786# vss nfet$276
Xnfet$269_0 m1_n8625_26174# vss m1_n8055_24542# vss nfet$269
Xnfet$262_7 m1_n7401_15478# m1_n7401_15478# m1_n927_19404# m1_n927_19404# m1_n695_20470#
+ vss nfet$262
Xnfet$255_6 m1_354_22513# m1_354_22513# m1_31535_22102# m1_31535_22102# m1_31771_21430#
+ vss nfet$255
Xnfet$253_3 m1_326_24346# m1_326_24346# vss vss m1_n192_24542# vss nfet$253
Xnfet$246_2 m1_12805_21786# vss m1_12935_21590# vss nfet$246
Xpfet$238_3 vdd vdd m1_34843_21786# m1_34093_19792# pfet$238
Xpfet$245_4 vdd vdd m1_26217_17714# m1_26676_16080# pfet$245
Xpfet$252_5 vdd m1_n6839_21786# vdd m1_n5764_21786# pfet$252
Xnfet$261_18 m1_23930_15778# m1_23930_15778# m1_23820_18030# m1_23820_18030# m1_24056_17358#
+ vss nfet$261
Xnfet$245_19 m1_n7513_20152# vss m1_1578_16080# vss nfet$245
Xnfet$251_0 m1_n1134_25662# m1_n910_23922# m1_n646_24542# vss nfet$251
Xpfet$236_0 vdd vdd m1_n646_24542# m1_n290_24224# pfet$236
Xpfet$233_14 vdd vdd m1_23486_19550# m1_21564_17714# pfet$233
Xpfet$228_69 vdd vdd m1_20721_15778# m1_17851_17714# pfet$228
Xpfet$228_14 vdd vdd m1_2092_17836# m1_1933_17343# pfet$228
Xpfet$228_25 vdd vdd m1_1709_17518# m1_1119_17714# pfet$228
Xpfet$228_36 vdd vdd m1_6116_17343# m1_9015_17714# pfet$228
Xpfet$228_47 vdd m1_11738_16080# m1_11271_18030# m1_10299_17343# pfet$228
Xpfet$228_58 vdd vdd m1_n3534_17714# m1_n3064_17714# pfet$228
Xpfet$230_26 vdd m1_n1927_20274# m1_n1927_20274# m1_17526_19550# m1_13198_17714# m1_13198_17714#
+ pfet$230
Xpfet$230_15 vdd vdd vdd m1_n59_19550# m1_n7401_15478# m1_n7401_15478# pfet$230
Xnfet$269_1 m1_n8625_26174# vss m1_n7082_23622# vss nfet$269
Xnfet$255_7 m1_3871_22513# m1_3871_22513# vss vss m1_31771_21430# vss nfet$255
Xnfet$262_8 m1_26063_15478# m1_26063_15478# m1_n3822_20130# m1_n3822_20130# m1_27441_20470#
+ vss nfet$262
Xnfet$253_4 m1_33174_24224# m1_33174_24224# m1_32818_24542# m1_32818_24542# m1_33272_24542#
+ vss nfet$253
Xnfet$246_3 m1_9288_21786# vss m1_9418_21590# vss nfet$246
Xpfet$238_4 vdd m1_34093_19792# vdd m1_32818_20470# pfet$238
Xpfet$245_5 vdd m1_26217_17714# vdd m1_27292_16202# pfet$245
Xpfet$252_6 vdd vdd m1_n6973_21481# m1_n6839_21786# pfet$252
Xnfet$244_0 m1_n3534_17714# m1_n3534_17714# vss vss m1_3454_20470# vss nfet$244
Xnfet$251_1 m1_n1271_25858# m1_n647_25662# m1_n910_23922# vss nfet$251
Xnfet$261_19 m1_23109_16202# m1_23109_16202# vss vss m1_22591_16398# vss nfet$261
Xpfet$236_1 vdd m1_n789_25858# vdd m1_814_25658# pfet$236
Xpfet$229_0 vdd vdd vdd m1_n674_22102# m1_n1133_21590# m1_n1133_21590# pfet$229
Xpfet$233_15 vdd vdd m1_22205_20152# m1_17697_15478# pfet$233
Xpfet$228_15 vdd vdd m1_5302_17714# m1_5761_16080# pfet$228
Xpfet$228_26 vdd vdd m1_4832_17714# m1_5302_17714# pfet$228
Xpfet$228_37 vdd m1_7555_16080# m1_7088_18030# m1_6116_17343# pfet$228
Xpfet$228_48 vdd vdd m1_n3064_17714# m1_n2605_16080# pfet$228
Xpfet$228_59 vdd vdd m1_n2605_16080# m1_n7513_20152# pfet$228
Xpfet$230_27 vdd vdd vdd m1_20407_19850# m1_22205_20152# m1_22205_20152# pfet$230
Xpfet$230_16 vdd vdd vdd m1_28077_19550# m1_26063_15478# m1_26063_15478# pfet$230
Xnfet$269_2 vss vss m1_n9336_24346# vss nfet$269
Xnfet$262_9 m1_29239_20152# m1_29239_20152# m1_n3822_20130# m1_n3822_20130# m1_28073_20470#
+ vss nfet$262
Xpfet$259_0 vdd vdd m1_n8145_21908# m1_n6839_20152# pfet$259
Xnfet$274_0 m1_n4485_21904# m1_n5764_21786# vss vss nfet$274
Xnfet$253_5 m1_33790_24346# m1_33790_24346# vss vss m1_33272_24542# vss nfet$253
Xpfet$245_6 vdd vdd m1_28003_18030# m1_28113_15778# pfet$245
Xpfet$238_5 vdd vdd m1_34093_19792# m1_32818_21586# pfet$238
Xpfet$252_7 vdd vdd m1_n6839_21786# m1_n6380_21786# pfet$252
Xnfet$246_4 m1_7522_21786# vss m1_8154_21786# vss nfet$246
Xnfet$244_1 m1_2384_19550# m1_2384_19550# vss vss m1_2822_20470# vss nfet$244
Xnfet$251_2 m1_n1271_25858# m1_814_25658# m1_1607_24542# vss nfet$251
Xpfet$236_2 vdd vdd m1_n789_25858# m1_326_24346# pfet$236
Xpfet$229_1 vdd m1_7388_22513# m1_7388_22513# m1_6988_22402# m1_7522_21786# m1_7522_21786#
+ pfet$229
Xpfet$233_16 vdd vdd m1_19969_19550# m1_17381_17714# pfet$233
Xpfet$241_0 vdd m1_34093_22102# vdd m1_28490_22513# pfet$241
Xpfet$228_16 vdd vdd m1_3989_15778# m1_1119_17714# pfet$228
Xpfet$228_27 vdd m1_2194_16202# m1_1709_17518# m1_2092_17836# pfet$228
Xpfet$228_38 vdd vdd m1_7088_18030# m1_7198_15778# pfet$228
Xpfet$228_49 vdd m1_n194_15778# m1_n811_16080# m1_n2091_17836# pfet$228
Xpfet$230_28 vdd vdd vdd m1_21043_19550# m1_17697_15478# m1_17697_15478# pfet$230
Xpfet$230_17 vdd m1_n3822_20130# m1_n3822_20130# m1_28077_19550# m1_25747_17714# m1_25747_17714#
+ pfet$230
Xnfet$269_3 fin vss m1_n10933_25858# vss nfet$269
Xnfet$243_10 m1_19839_21786# m1_19839_21786# m1_21456_22513# m1_21456_22513# m1_21060_21586#
+ vss nfet$243
Xnfet$274_1 m1_n5227_21418# vss m1_n5764_21786# vss nfet$274
Xnfet$267_0 m1_n7082_23622# m1_n6856_24542# vss vss nfet$267
Xnfet$253_6 m1_33790_24346# m1_33790_24346# m1_32675_25947# m1_32675_25947# m1_34737_25502#
+ vss nfet$253
Xpfet$245_7 vdd m1_28003_18030# vdd m1_26676_16080# pfet$245
Xnfet$246_5 m1_488_21786# vss m1_1120_21786# vss nfet$246
Xpfet$238_6 vdd vdd m1_31535_19792# m1_14422_22513# pfet$238
Xnfet$251_3 m1_n1134_25662# m1_n290_24224# m1_814_25658# vss nfet$251
Xpfet$236_3 vdd m1_n646_24542# vdd m1_326_24346# pfet$236
Xnfet$244_2 m1_5901_19550# m1_5901_19550# vss vss m1_6339_20470# vss nfet$244
Xpfet$229_2 vdd m1_7388_22513# m1_7388_22513# m1_6360_22102# m1_8154_21786# m1_8154_21786#
+ pfet$229
Xpfet$233_17 vdd vdd m1_25722_20152# m1_21880_15478# pfet$233
Xpfet$241_1 vdd vdd m1_34093_22102# m1_34843_21786# pfet$241
Xnfet$246_10 m1_21590_21786# vss m1_22222_21786# vss nfet$246
Xpfet$234_0 vdd vdd m1_n7401_15478# sd9 pfet$234
Xpfet$228_17 vdd vdd m1_n2091_17836# m1_n2250_17343# pfet$228
Xpfet$228_28 vdd m1_2905_18030# vdd m1_1578_16080# pfet$228
Xpfet$228_39 vdd m1_7088_18030# vdd m1_5761_16080# pfet$228
Xpfet$230_29 vdd vdd vdd m1_23924_19850# m1_25722_20152# m1_25722_20152# pfet$230
Xpfet$230_18 vdd vdd vdd m1_27441_19850# m1_29239_20152# m1_29239_20152# pfet$230
Xnfet$269_4 m1_n10572_23922# vss m1_n9952_24224# vss nfet$269
Xnfet$243_11 m1_19969_21590# m1_19969_21590# m1_21456_22513# m1_21456_22513# m1_20428_21586#
+ vss nfet$243
Xnfet$274_2 m1_n6839_21786# vss m1_n6973_21481# vss nfet$274
Xnfet$267_1 m1_n8283_19850# vss m1_n6856_24542# vss nfet$267
Xnfet$254_10 m1_21590_21786# m1_21590_21786# vss vss m1_20428_21586# vss nfet$254
Xnfet$253_7 m1_34278_25658# m1_34278_25658# vss vss m1_34737_25502# vss nfet$253
Xnfet$246_6 m1_5771_21786# vss m1_5901_21590# vss nfet$246
Xpfet$238_7 vdd vdd m1_31535_22102# m1_354_22513# pfet$238
Xnfet$249_10 m1_26217_17714# vss m1_29087_15778# vss nfet$249
Xpfet$236_4 vdd vdd m1_32675_25947# m1_33790_24346# pfet$236
Xnfet$251_4 m1_32193_25858# m1_34278_25658# m1_35071_24542# vss nfet$251
Xnfet$244_3 m1_4832_17714# m1_4832_17714# vss vss m1_10488_20470# vss nfet$244
Xpfet$229_3 vdd m1_9645_21447# m1_9645_21447# m1_10505_22402# m1_11039_21786# m1_11039_21786#
+ pfet$229
Xnfet$242_0 m1_3394_25858# vss m1_5790_24542# vss nfet$242
Xpfet$241_2 vdd vdd m1_30256_22102# m1_7388_22513# pfet$241
Xnfet$246_11 m1_18073_21786# vss m1_18705_21786# vss nfet$246
Xpfet$234_1 vdd vdd m1_21880_15478# sd2 pfet$234
Xpfet$227_0 vdd vdd m1_3049_25662# m1_2912_25858# pfet$227
Xnfet$262_10 m1_9331_15478# m1_9331_15478# m1_n3822_21786# m1_n3822_21786# m1_13373_20470#
+ vss nfet$262
Xpfet$228_18 vdd m1_1119_17714# vdd m1_2194_16202# pfet$228
Xpfet$228_29 vdd vdd m1_1578_16080# m1_n7513_20152# pfet$228
Xpfet$230_19 vdd m1_n3822_20130# m1_n3822_20130# m1_27441_19850# m1_27003_19550# m1_27003_19550#
+ pfet$230
Xnfet$269_5 m1_n10933_25858# vss m1_n10796_25662# vss nfet$269
Xnfet$243_12 m1_16322_21786# m1_16322_21786# m1_17939_22513# m1_17939_22513# m1_17543_21586#
+ vss nfet$243
Xnfet$254_11 m1_22222_21786# m1_22222_21786# vss vss m1_21060_21586# vss nfet$254
Xnfet$246_7 m1_4005_21786# vss m1_4637_21786# vss nfet$246
Xnfet$272_0 m1_n7186_25858# vss m1_n7320_25516# vss nfet$272
Xnfet$249_11 m1_27031_17343# vss m1_27190_17836# vss nfet$249
Xpfet$257_0 vdd vdd m1_n5227_20152# m1_n2543_20130# pfet$257
Xnfet$251_5 m1_32330_25662# m1_33174_24224# m1_34278_25658# vss nfet$251
Xnfet$244_4 m1_9418_19550# m1_9418_19550# vss vss m1_9856_20470# vss nfet$244
Xpfet$236_5 vdd m1_32675_25947# vdd m1_34278_25658# pfet$236
Xpfet$229_4 vdd vdd vdd m1_9877_22102# m1_9418_21590# m1_9418_21590# pfet$229
Xpfet$234_2 vdd vdd m1_26063_15478# sd1 pfet$234
Xpfet$241_3 vdd m1_31535_22102# vdd m1_3871_22513# pfet$241
Xpfet$227_1 vdd m1_3536_25662# m1_3273_23922# m1_3049_25662# pfet$227
Xnfet$242_1 m1_2912_25858# m1_4997_25658# m1_5790_24542# vss nfet$242
Xnfet$246_12 m1_14556_21786# vss m1_15188_21786# vss nfet$246
Xnfet$262_11 m1_15171_20152# m1_15171_20152# m1_n3822_21786# m1_n3822_21786# m1_14005_20470#
+ vss nfet$262
Xpfet$228_19 vdd m1_3015_15778# m1_2194_16202# m1_1933_17343# pfet$228
Xnfet$269_6 m1_n10452_25858# vss m1_n10309_25662# vss nfet$269
Xnfet$243_13 m1_16452_21590# m1_16452_21590# m1_17939_22513# m1_17939_22513# m1_16911_21586#
+ vss nfet$243
Xnfet$254_12 m1_18073_21786# m1_18073_21786# vss vss m1_16911_21586# vss nfet$254
Xnfet$246_8 m1_2254_21786# vss m1_2384_21590# vss nfet$246
Xnfet$265_0 m1_n5351_15778# m1_n5351_15778# m1_n5461_18030# m1_n5461_18030# m1_n5225_17358#
+ vss nfet$265
Xnfet$272_1 m1_n6856_24542# vss m1_n6111_25858# vss nfet$272
Xnfet$249_12 m1_28470_16080# vss m1_28113_15778# vss nfet$249
Xpfet$257_1 vdd m1_n4485_20152# vdd m1_n3206_20274# pfet$257
Xnfet$251_6 m1_32193_25858# m1_32817_25662# m1_32554_23922# vss nfet$251
Xnfet$244_5 m1_649_17714# m1_649_17714# vss vss m1_6971_20470# vss nfet$244
Xpfet$236_6 vdd vdd m1_32818_24542# m1_33174_24224# pfet$236
Xpfet$229_5 vdd m1_9645_21447# m1_9645_21447# m1_9877_22102# m1_11671_21786# m1_11671_21786#
+ pfet$229
Xpfet$241_4 vdd m1_30256_22102# vdd m1_9645_21447# pfet$241
Xnfet$242_2 m1_n7513_20152# vss m1_4509_24346# vss nfet$242
Xnfet$246_13 m1_16322_21786# vss m1_16452_21590# vss nfet$246
Xnfet$262_12 m1_18688_20152# m1_18688_20152# m1_n1927_20274# m1_n1927_20274# m1_17522_20470#
+ vss nfet$262
Xpfet$227_2 vdd vdd m1_3394_25858# m1_4509_24346# pfet$227
Xpfet$232_0 vdd vdd m1_n6274_17836# m1_n6433_17343# pfet$232
Xnfet$269_7 m1_n7320_25516# vss m1_n2567_23922# vss nfet$269
Xpfet$229_30 vdd vdd vdd m1_17539_22402# m1_16322_21786# m1_16322_21786# pfet$229
Xnfet$243_14 m1_12805_21786# m1_12805_21786# m1_14422_22513# m1_14422_22513# m1_14026_21586#
+ vss nfet$243
Xnfet$254_13 m1_18705_21786# m1_18705_21786# vss vss m1_17543_21586# vss nfet$254
Xnfet$246_9 m1_23356_21786# vss m1_23486_21590# vss nfet$246
Xnfet$258_0 m1_34093_19792# vss m1_34843_21786# vss nfet$258
Xnfet$265_1 m1_n6788_16080# m1_n6788_16080# vss vss m1_n5225_17358# vss nfet$265
Xnfet$249_13 m1_26217_17714# vss m1_25747_17714# vss nfet$249
Xpfet$257_2 vdd m1_n5227_20152# vdd m1_n1927_20274# pfet$257
Xnfet$251_7 m1_32330_25662# m1_32554_23922# m1_32818_24542# vss nfet$251
Xnfet$244_6 m1_n1133_19550# m1_n1133_19550# vss vss m1_n695_20470# vss nfet$244
Xpfet$236_7 vdd m1_32818_24542# vdd m1_33790_24346# pfet$236
Xpfet$229_6 vdd vdd vdd m1_10505_22402# m1_9288_21786# m1_9288_21786# pfet$229
Xnfet$242_3 m1_488_21786# vss m1_2912_25858# vss nfet$242
Xnfet$246_14 m1_19839_21786# vss m1_19969_21590# vss nfet$246
Xnfet$262_13 m1_13514_15478# m1_13514_15478# m1_n1927_20274# m1_n1927_20274# m1_16890_20470#
+ vss nfet$262
Xpfet$227_3 vdd m1_3394_25858# vdd m1_4997_25658# pfet$227
Xpfet$232_1 vdd vdd m1_n4377_15778# m1_n7247_17714# pfet$232
Xnfet$269_8 m1_n4623_25487# vss m1_n4464_25980# vss nfet$269
Xpfet$229_31 vdd vdd vdd m1_27462_22102# m1_27003_21590# m1_27003_21590# pfet$229
Xpfet$229_20 vdd vdd vdd m1_20428_22102# m1_19969_21590# m1_19969_21590# pfet$229
Xnfet$243_15 m1_26873_21786# m1_26873_21786# m1_28490_22513# m1_28490_22513# m1_28094_21586#
+ vss nfet$243
Xpfet$231_10 vdd vdd m1_23486_21590# m1_23356_21786# pfet$231
Xnfet$254_14 m1_15188_21786# m1_15188_21786# vss vss m1_14026_21586# vss nfet$254
Xnfet$258_1 m1_30256_19792# vss m1_32818_20470# vss nfet$258
Xnfet$265_2 m1_n6788_16080# m1_n6788_16080# m1_n7247_17714# m1_n7247_17714# m1_n6690_16398#
+ vss nfet$265
Xpfet$257_3 vdd m1_n6839_20152# vdd m1_n927_19404# pfet$257
Xnfet$244_7 m1_n7383_17599# m1_n7383_17599# vss vss m1_n63_20470# vss nfet$244
Xnfet$270_0 m1_n9952_24224# m1_n9952_24224# m1_n10308_24542# m1_n10308_24542# m1_n9854_24542#
+ vss nfet$270
Xpfet$229_7 vdd m1_354_22513# m1_354_22513# m1_n674_22102# m1_1120_21786# m1_1120_21786#
+ pfet$229
Xpfet$255_0 vdd vdd vdd m1_n8047_19550# m1_n7513_20152# m1_n7513_20152# pfet$255
Xnfet$242_4 m1_2912_25858# vss m1_3049_25662# vss nfet$242
Xnfet$246_15 m1_28624_21786# vss m1_29256_21786# vss nfet$246
Xnfet$262_14 m1_22205_20152# m1_22205_20152# m1_n2543_20130# m1_n2543_20130# m1_21039_20470#
+ vss nfet$262
Xpfet$227_4 vdd vdd m1_3893_24224# m1_3273_23922# pfet$227
Xpfet$232_2 vdd vdd m1_n5351_15778# m1_n4994_16080# pfet$232
Xnfet$269_9 m1_n3184_24224# vss m1_n3541_23922# vss nfet$269
Xpfet$229_32 vdd m1_28490_22513# m1_28490_22513# m1_28090_22402# m1_28624_21786# m1_28624_21786#
+ pfet$229
Xpfet$229_21 vdd vdd vdd m1_21056_22402# m1_19839_21786# m1_19839_21786# pfet$229
Xpfet$229_10 vdd m1_3871_22513# m1_3871_22513# m1_2843_22102# m1_4637_21786# m1_4637_21786#
+ pfet$229
Xnfet$243_16 m1_27003_21590# m1_27003_21590# m1_28490_22513# m1_28490_22513# m1_27462_21586#
+ vss nfet$243
Xpfet$231_11 vdd vdd m1_18705_21786# m1_18073_21786# pfet$231
Xnfet$254_15 m1_14556_21786# m1_14556_21786# vss vss m1_13394_21586# vss nfet$254
Xnfet$258_2 m1_31535_19792# m1_32818_20470# vss vss nfet$258
Xnfet$265_3 m1_n6172_16202# m1_n6172_16202# vss vss m1_n6690_16398# vss nfet$265
Xpfet$257_4 vdd vdd m1_n6839_20152# m1_n6973_21481# pfet$257
Xnfet$263_0 m1_35837_22102# vss m1_n7513_20152# vss nfet$263
Xnfet$244_8 m1_27003_19550# m1_27003_19550# vss vss m1_27441_20470# vss nfet$244
Xnfet$270_1 m1_n9336_24346# m1_n9336_24346# m1_n8625_26174# m1_n8625_26174# m1_n8389_25502#
+ vss nfet$270
Xpfet$229_8 vdd vdd vdd m1_6360_22102# m1_5901_21590# m1_5901_21590# pfet$229
Xpfet$255_1 vdd m1_n8283_19850# m1_n8283_19850# m1_n8047_19550# m1_n8283_20611# m1_n8283_20611#
+ pfet$255
Xpfet$248_0 vdd vdd vdd m1_n6624_23622# m1_n7082_23622# m1_n7082_23622# pfet$248
Xnfet$242_5 m1_2912_25858# m1_3536_25662# m1_3273_23922# vss nfet$242
Xnfet$246_16 m1_26873_21786# vss m1_27003_21590# vss nfet$246
Xpfet$227_5 vdd m1_3893_24224# m1_4997_25658# m1_2912_25858# pfet$227
Xnfet$262_15 m1_17697_15478# m1_17697_15478# m1_n2543_20130# m1_n2543_20130# m1_20407_20470#
+ vss nfet$262
Xpfet$232_3 vdd vdd m1_n6657_17518# m1_n7247_17714# pfet$232
Xpfet$228_110 vdd vdd m1_10458_17836# m1_10299_17343# pfet$228
Xpfet$229_33 vdd m1_28490_22513# m1_28490_22513# m1_27462_22102# m1_29256_21786# m1_29256_21786#
+ pfet$229
Xpfet$229_22 vdd m1_21456_22513# m1_21456_22513# m1_20428_22102# m1_22222_21786# m1_22222_21786#
+ pfet$229
Xpfet$229_11 vdd vdd vdd m1_2843_22102# m1_2384_21590# m1_2384_21590# pfet$229
Xnfet$243_17 m1_12935_21590# m1_12935_21590# m1_14422_22513# m1_14422_22513# m1_13394_21586#
+ vss nfet$243
Xpfet$230_0 vdd m1_2590_19404# m1_2590_19404# m1_3458_19550# m1_n3534_17714# m1_n3534_17714#
+ pfet$230
Xpfet$231_12 vdd vdd m1_16452_21590# m1_16322_21786# pfet$231
Xnfet$254_16 m1_28624_21786# m1_28624_21786# vss vss m1_27462_21586# vss nfet$254
Xnfet$258_3 m1_30256_22102# vss m1_32818_21586# vss nfet$258
Xnfet$265_4 m1_28113_15778# m1_28113_15778# m1_28003_18030# m1_28003_18030# m1_28239_17358#
+ vss nfet$265
Xnfet$244_9 m1_25747_17714# m1_25747_17714# vss vss m1_28073_20470# vss nfet$244
Xnfet$256_0 m1_34843_21786# m1_34843_21786# m1_34093_22102# m1_34093_22102# m1_34329_21430#
+ vss nfet$256
Xpfet$255_2 vdd m1_n8283_20611# m1_n8283_20611# m1_n8047_22344# m1_n8145_21908# m1_n8145_21908#
+ pfet$255
Xnfet$270_2 m1_n8848_25658# m1_n8848_25658# vss vss m1_n8389_25502# vss nfet$270
Xpfet$253_10 vdd vdd m1_n10933_25858# fin pfet$253
Xpfet$248_1 vdd m1_n6856_24542# m1_n6856_24542# m1_n6624_23622# m1_n8283_19850# m1_n8283_19850#
+ pfet$248
Xpfet$229_9 vdd m1_3871_22513# m1_3871_22513# m1_3471_22402# m1_4005_21786# m1_4005_21786#
+ pfet$229
Xpfet$227_6 vdd vdd m1_3536_25662# m1_3394_25858# pfet$227
Xnfet$242_6 m1_3049_25662# m1_3893_24224# m1_4997_25658# vss nfet$242
Xnfet$246_17 m1_25107_21786# vss m1_25739_21786# vss nfet$246
Xnfet$262_16 m1_25722_20152# m1_25722_20152# m1_n3206_20274# m1_n3206_20274# m1_24556_20470#
+ vss nfet$262
Xpfet$232_4 vdd vdd m1_n6433_17343# m1_n3534_17714# pfet$232
Xpfet$229_12 vdd vdd vdd m1_3471_22402# m1_2254_21786# m1_2254_21786# pfet$229
Xpfet$229_34 vdd vdd vdd m1_28090_22402# m1_26873_21786# m1_26873_21786# pfet$229
Xpfet$229_23 vdd vdd vdd m1_23945_22102# m1_23486_21590# m1_23486_21590# pfet$229
Xpfet$228_100 vdd vdd m1_23820_18030# m1_23930_15778# pfet$228
Xpfet$230_1 vdd vdd vdd m1_2822_19850# m1_4620_20152# m1_4620_20152# pfet$230
Xpfet$231_13 vdd vdd m1_15188_21786# m1_14556_21786# pfet$231
Xnfet$254_17 m1_29256_21786# m1_29256_21786# vss vss m1_28094_21586# vss nfet$254
Xnfet$265_5 m1_26676_16080# m1_26676_16080# vss vss m1_28239_17358# vss nfet$265
Xnfet$256_1 m1_28490_22513# m1_28490_22513# vss vss m1_34329_21430# vss nfet$256
Xnfet$249_0 m1_n3534_17714# vss m1_n6433_17343# vss nfet$249
Xnfet$270_3 m1_n9336_24346# m1_n9336_24346# vss vss m1_n9854_24542# vss nfet$270
Xpfet$253_11 vdd vdd m1_n9336_24346# vss pfet$253
Xpfet$255_3 vdd vdd vdd m1_n8047_22344# m1_n8283_19850# m1_n8283_19850# pfet$255
Xnfet$242_7 m1_3049_25662# m1_3273_23922# m1_3537_24542# vss nfet$242
Xnfet$262_17 m1_21880_15478# m1_21880_15478# m1_n3206_20274# m1_n3206_20274# m1_23924_20470#
+ vss nfet$262
Xpfet$227_7 vdd vdd m1_7232_25662# m1_7095_25858# pfet$227
Xpfet$253_0 vdd vdd m1_n10796_25662# m1_n10933_25858# pfet$253
Xpfet$232_5 vdd vdd m1_n6788_16080# m1_n7513_20152# pfet$232
Xpfet$229_35 vdd vdd vdd m1_13394_22102# m1_12935_21590# m1_12935_21590# pfet$229
Xpfet$229_24 vdd m1_17939_22513# m1_17939_22513# m1_16911_22102# m1_18705_21786# m1_18705_21786#
+ pfet$229
Xpfet$228_101 vdd vdd m1_19637_18030# m1_19747_15778# pfet$228
Xpfet$229_13 vdd vdd vdd m1_6988_22402# m1_5771_21786# m1_5771_21786# pfet$229
Xpfet$230_2 vdd m1_2590_19404# m1_2590_19404# m1_2822_19850# m1_2384_19550# m1_2384_19550#
+ pfet$230
Xpfet$231_14 vdd vdd m1_19969_21590# m1_19839_21786# pfet$231
Xnfet$265_6 m1_27292_16202# m1_27292_16202# vss vss m1_26774_16398# vss nfet$265
Xnfet$256_2 m1_9645_21447# m1_9645_21447# vss vss m1_30492_21430# vss nfet$256
Xnfet$249_1 m1_n7513_20152# vss m1_n6788_16080# vss nfet$249
Xnfet$270_4 m1_n4978_24224# m1_n4978_24224# m1_n10452_25858# m1_n10452_25858# m1_n4880_24542#
+ vss nfet$270
Xpfet$253_12 vdd vdd m1_n7082_23622# m1_n8625_26174# pfet$253
Xpfet$227_90 vdd vdd m1_24309_25858# m1_25424_24346# pfet$227
Xnfet$242_8 m1_3394_25858# vss m1_3536_25662# vss nfet$242
Xpfet$227_8 vdd vdd m1_8076_24224# m1_7456_23922# pfet$227
Xnfet$261_0 m1_7198_15778# m1_7198_15778# m1_7088_18030# m1_7088_18030# m1_7324_17358#
+ vss nfet$261
Xpfet$246_0 vdd m1_n4377_15778# m1_n4994_16080# m1_n6274_17836# pfet$246
Xpfet$253_1 vdd vdd m1_n10309_25662# m1_n10452_25858# pfet$253
Xpfet$232_6 vdd vdd m1_n7383_17599# m1_n7247_17714# pfet$232
Xpfet$229_25 vdd m1_17939_22513# m1_17939_22513# m1_17539_22402# m1_18073_21786# m1_18073_21786#
+ pfet$229
Xpfet$228_102 vdd vdd m1_13198_17714# m1_13668_17714# pfet$228
Xpfet$229_14 vdd vdd vdd m1_n46_22402# m1_n1263_21786# m1_n1263_21786# pfet$229
Xpfet$230_3 vdd vdd vdd m1_3458_19550# m1_n3218_15478# m1_n3218_15478# pfet$230
Xpfet$231_15 vdd vdd m1_27003_21590# m1_26873_21786# pfet$231
Xnfet$265_7 m1_26676_16080# m1_26676_16080# m1_26217_17714# m1_26217_17714# m1_26774_16398#
+ vss nfet$265
Xnfet$256_3 m1_7388_22513# m1_7388_22513# m1_30256_22102# m1_30256_22102# m1_30492_21430#
+ vss nfet$256
Xnfet$249_2 m1_n4994_16080# vss m1_n5351_15778# vss nfet$249
Xnfet$270_5 m1_n4362_24346# m1_n4362_24346# vss vss m1_n4880_24542# vss nfet$270
Xpfet$253_13 vdd vdd m1_n8055_24542# m1_n8625_26174# pfet$253
Xpfet$227_91 vdd vdd m1_23356_21786# pd8 pfet$227
Xpfet$227_80 vdd vdd m1_17058_24346# m1_n7513_20152# pfet$227
Xnfet$241_20 m1_21241_24346# m1_21241_24346# m1_20126_25858# m1_20126_25858# m1_22188_25502#
+ vss nfet$241
Xnfet$242_9 m1_3273_23922# vss m1_3893_24224# vss nfet$242
Xpfet$227_9 vdd m1_7719_25662# m1_7456_23922# m1_7232_25662# pfet$227
Xnfet$261_1 m1_5761_16080# m1_5761_16080# vss vss m1_7324_17358# vss nfet$261
Xnfet$254_0 m1_11039_21786# m1_11039_21786# vss vss m1_9877_21586# vss nfet$254
Xpfet$246_1 vdd m1_n5351_15778# m1_n6172_16202# m1_n6433_17343# pfet$246
Xpfet$253_2 vdd vdd m1_n9952_24224# m1_n10572_23922# pfet$253
Xpfet$239_0 vdd m1_n647_25662# m1_n910_23922# m1_n1134_25662# pfet$239
Xpfet$232_7 vdd vdd m1_27190_17836# m1_27031_17343# pfet$232
Xpfet$229_26 vdd vdd vdd m1_16911_22102# m1_16452_21590# m1_16452_21590# pfet$229
Xpfet$228_103 vdd m1_14743_16202# m1_14258_17518# m1_14641_17836# pfet$228
Xpfet$229_15 vdd m1_354_22513# m1_354_22513# m1_n46_22402# m1_488_21786# m1_488_21786#
+ pfet$229
Xpfet$230_4 vdd m1_6107_19404# m1_6107_19404# m1_6339_19850# m1_5901_19550# m1_5901_19550#
+ pfet$230
Xpfet$231_16 vdd vdd m1_29256_21786# m1_28624_21786# pfet$231
Xnfet$270_6 m1_n4978_24224# m1_n4978_24224# vss vss m1_n3415_25502# vss nfet$270
Xpfet$227_92 vdd vdd m1_28492_25858# m1_29607_24346# pfet$227
Xpfet$227_81 vdd vdd m1_18339_24542# m1_15943_25858# pfet$227
Xpfet$227_70 vdd vdd m1_14156_24542# m1_11760_25858# pfet$227
Xnfet$249_3 m1_n6433_17343# vss m1_n6274_17836# vss nfet$249
Xnfet$241_21 m1_28991_24224# m1_28991_24224# m1_28635_24542# m1_28635_24542# m1_29089_24542#
+ vss nfet$241
Xnfet$241_10 m1_17546_25658# m1_17546_25658# vss vss m1_18005_25502# vss nfet$241
Xnfet$247_0 m1_n3534_17714# vss m1_2384_19550# vss nfet$247
Xnfet$261_2 m1_9944_16080# m1_9944_16080# vss vss m1_11507_17358# vss nfet$261
Xnfet$254_1 m1_11671_21786# m1_11671_21786# vss vss m1_10509_21586# vss nfet$254
Xpfet$246_2 vdd m1_n4994_16080# m1_n5461_18030# m1_n6433_17343# pfet$246
Xpfet$253_3 vdd vdd m1_n4978_24224# vss pfet$253
Xpfet$239_1 vdd m1_n910_23922# m1_n646_24542# m1_n1271_25858# pfet$239
Xpfet$232_8 vdd vdd m1_28113_15778# m1_28470_16080# pfet$232
Xpfet$251_0 vdd vdd m1_n8625_26174# m1_n9336_24346# pfet$251
Xpfet$229_27 vdd m1_14422_22513# m1_14422_22513# m1_14022_22402# m1_14556_21786# m1_14556_21786#
+ pfet$229
Xpfet$229_16 vdd m1_24973_22513# m1_24973_22513# m1_23945_22102# m1_25739_21786# m1_25739_21786#
+ pfet$229
Xpfet$228_104 vdd vdd m1_14127_16080# m1_n7513_20152# pfet$228
Xpfet$230_5 vdd vdd vdd m1_n695_19850# m1_1103_20152# m1_1103_20152# pfet$230
Xpfet$231_17 vdd vdd m1_25739_21786# m1_25107_21786# pfet$231
Xnfet$244_10 m1_9015_17714# m1_9015_17714# vss vss m1_14005_20470# vss nfet$244
Xnfet$277_0 m1_n6839_20152# vss m1_n8145_21908# vss nfet$277
Xnfet$249_4 m1_n7247_17714# vss m1_n4377_15778# vss nfet$249
Xnfet$270_7 m1_n3541_23922# m1_n3541_23922# m1_n3651_26174# m1_n3651_26174# m1_n3415_25502#
+ vss nfet$270
Xnfet$241_22 m1_29607_24346# m1_29607_24346# vss vss m1_29089_24542# vss nfet$241
Xpfet$227_93 vdd m1_28991_24224# m1_30095_25658# m1_28010_25858# pfet$227
Xpfet$227_82 vdd vdd m1_21241_24346# m1_n7513_20152# pfet$227
Xpfet$227_71 vdd vdd m1_11039_21786# m1_11760_25858# pfet$227
Xpfet$227_60 vdd vdd m1_20126_25858# m1_21241_24346# pfet$227
Xnfet$241_11 m1_16442_24224# m1_16442_24224# m1_16086_24542# m1_16086_24542# m1_16540_24542#
+ vss nfet$241
Xnfet$247_1 m1_n3218_15478# vss m1_4620_20152# vss nfet$247
Xnfet$261_3 m1_11381_15778# m1_11381_15778# m1_11271_18030# m1_11271_18030# m1_11507_17358#
+ vss nfet$261
Xnfet$254_2 m1_8154_21786# m1_8154_21786# vss vss m1_6992_21586# vss nfet$254
Xpfet$246_3 vdd m1_n6172_16202# m1_n6657_17518# m1_n6274_17836# pfet$246
Xpfet$253_4 vdd vdd m1_n5571_25662# m1_n10452_25858# pfet$253
Xpfet$239_2 vdd m1_n290_24224# m1_814_25658# m1_n1271_25858# pfet$239
Xpfet$232_9 vdd vdd m1_29087_15778# m1_26217_17714# pfet$232
Xpfet$229_28 vdd m1_14422_22513# m1_14422_22513# m1_13394_22102# m1_15188_21786# m1_15188_21786#
+ pfet$229
Xpfet$229_17 vdd m1_21456_22513# m1_21456_22513# m1_21056_22402# m1_21590_21786# m1_21590_21786#
+ pfet$229
Xpfet$244_0 vdd m1_32818_20470# m1_32818_20470# m1_33050_19550# m1_30256_19792# m1_30256_19792#
+ pfet$244
Xnfet$247_10 m1_26063_15478# vss m1_29239_20152# vss nfet$247
Xpfet$251_1 vdd m1_n8625_26174# vdd m1_n8848_25658# pfet$251
Xpfet$228_105 vdd vdd m1_14258_17518# m1_13668_17714# pfet$228
Xpfet$230_6 vdd vdd vdd m1_6339_19850# m1_8137_20152# m1_8137_20152# pfet$230
Xnfet$244_11 m1_13198_17714# m1_13198_17714# vss vss m1_17522_20470# vss nfet$244
Xnfet$249_5 m1_n7247_17714# vss m1_n6657_17518# vss nfet$249
Xnfet$241_23 m1_25424_24346# m1_25424_24346# m1_24309_25858# m1_24309_25858# m1_26371_25502#
+ vss nfet$241
Xpfet$227_94 vdd m1_28492_25858# vdd m1_30095_25658# pfet$227
Xpfet$227_83 vdd m1_21729_25658# m1_22522_24542# m1_19781_25662# pfet$227
Xpfet$227_72 vdd m1_13363_25658# m1_14156_24542# m1_11415_25662# pfet$227
Xpfet$227_61 vdd m1_24452_24542# vdd m1_25424_24346# pfet$227
Xpfet$227_50 vdd vdd m1_20268_25662# m1_20126_25858# pfet$227
Xnfet$241_12 m1_17058_24346# m1_17058_24346# m1_15943_25858# m1_15943_25858# m1_18005_25502#
+ vss nfet$241
Xnfet$261_4 m1_10560_16202# m1_10560_16202# vss vss m1_10042_16398# vss nfet$261
Xpfet$246_4 vdd m1_28113_15778# m1_27292_16202# m1_27031_17343# pfet$246
Xpfet$239_3 vdd m1_814_25658# m1_1607_24542# m1_n1134_25662# pfet$239
Xnfet$247_2 m1_n7401_15478# vss m1_1103_20152# vss nfet$247
Xpfet$253_5 vdd vdd m1_n4847_25662# m1_n10452_25858# pfet$253
Xnfet$254_3 m1_7522_21786# m1_7522_21786# vss vss m1_6360_21586# vss nfet$254
Xnfet$252_0 pd1 vss m1_n1263_21786# vss nfet$252
Xpfet$237_0 vdd vdd vdd m1_33050_22344# m1_31535_22102# m1_31535_22102# pfet$237
Xnfet$247_11 m1_9331_15478# vss m1_15171_20152# vss nfet$247
Xpfet$244_1 vdd vdd vdd m1_33050_19550# m1_31535_19792# m1_31535_19792# pfet$244
Xpfet$251_2 vdd m1_n3651_26174# vdd m1_n4978_24224# pfet$251
Xpfet$229_29 vdd vdd vdd m1_14022_22402# m1_12805_21786# m1_12805_21786# pfet$229
Xpfet$229_18 vdd vdd vdd m1_24573_22402# m1_23356_21786# m1_23356_21786# pfet$229
Xpfet$228_106 vdd vdd m1_14482_17343# m1_17381_17714# pfet$228
Xpfet$230_7 vdd vdd vdd m1_6975_19550# m1_965_15478# m1_965_15478# pfet$230
Xnfet$244_12 m1_16452_19550# m1_16452_19550# vss vss m1_16890_20470# vss nfet$244
Xnfet$249_6 m1_n7247_17714# vss m1_n7383_17599# vss nfet$249
Xpfet$227_95 vdd vdd m1_28991_24224# m1_28371_23922# pfet$227
Xpfet$227_84 vdd vdd m1_23827_25858# m1_18073_21786# pfet$227
Xpfet$227_73 vdd m1_16086_24542# vdd m1_17058_24346# pfet$227
Xpfet$227_62 vdd vdd m1_24452_24542# m1_24808_24224# pfet$227
Xpfet$227_51 vdd vdd m1_20625_24224# m1_20005_23922# pfet$227
Xpfet$227_40 vdd vdd m1_11760_25858# m1_12875_24346# pfet$227
Xnfet$241_24 m1_30095_25658# m1_30095_25658# vss vss m1_30554_25502# vss nfet$241
Xnfet$241_13 m1_13363_25658# m1_13363_25658# vss vss m1_13822_25502# vss nfet$241
Xpfet$246_5 vdd m1_29087_15778# m1_28470_16080# m1_27190_17836# pfet$246
Xnfet$247_3 m1_649_17714# vss m1_5901_19550# vss nfet$247
Xnfet$261_5 m1_9944_16080# m1_9944_16080# m1_9485_17714# m1_9485_17714# m1_10042_16398#
+ vss nfet$261
Xpfet$253_6 vdd vdd m1_n4623_25487# fin pfet$253
Xnfet$254_4 m1_1120_21786# m1_1120_21786# vss vss m1_n42_21586# vss nfet$254
Xpfet$239_4 vdd m1_33174_24224# m1_34278_25658# m1_32193_25858# pfet$239
Xnfet$252_1 pd2 vss m1_2254_21786# vss nfet$252
Xnfet$245_0 m1_9485_17714# vss m1_9015_17714# vss nfet$245
Xpfet$244_2 vdd m1_32818_21586# m1_32818_21586# m1_33050_22344# m1_30256_22102# m1_30256_22102#
+ pfet$244
Xnfet$247_12 m1_13514_15478# vss m1_18688_20152# vss nfet$247
Xpfet$251_3 vdd vdd m1_n3651_26174# m1_n3541_23922# pfet$251
Xpfet$229_19 vdd m1_24973_22513# m1_24973_22513# m1_24573_22402# m1_25107_21786# m1_25107_21786#
+ pfet$229
Xpfet$228_107 vdd m1_15921_16080# m1_15454_18030# m1_14482_17343# pfet$228
Xpfet$230_8 vdd m1_9624_19404# m1_9624_19404# m1_10492_19550# m1_4832_17714# m1_4832_17714#
+ pfet$230
Xnfet$244_13 m1_19969_19550# m1_19969_19550# vss vss m1_20407_20470# vss nfet$244
Xnfet$269_10 vss vss m1_n4978_24224# vss nfet$269
Xnfet$249_7 m1_26217_17714# vss m1_26807_17518# vss nfet$249
Xpfet$227_96 vdd m1_28635_24542# vdd m1_29607_24346# pfet$227
Xpfet$227_85 vdd m1_24188_23922# m1_24452_24542# m1_23827_25858# pfet$227
Xpfet$227_74 vdd vdd m1_14556_21786# m1_15943_25858# pfet$227
Xpfet$227_63 vdd vdd m1_19781_25662# m1_19644_25858# pfet$227
Xpfet$227_52 vdd m1_20268_25662# m1_20005_23922# m1_19781_25662# pfet$227
Xpfet$227_41 vdd vdd m1_9288_21786# pd4 pfet$227
Xpfet$227_30 vdd vdd m1_2912_25858# m1_488_21786# pfet$227
Xnfet$275_0 m1_n927_19404# m1_n927_19404# vss vss m1_n6282_20470# vss nfet$275
Xnfet$241_25 m1_29607_24346# m1_29607_24346# m1_28492_25858# m1_28492_25858# m1_30554_25502#
+ vss nfet$241
Xnfet$241_14 m1_12875_24346# m1_12875_24346# m1_11760_25858# m1_11760_25858# m1_13822_25502#
+ vss nfet$241
Xnfet$247_4 m1_4832_17714# vss m1_9418_19550# vss nfet$247
Xnfet$261_6 m1_1578_16080# m1_1578_16080# vss vss m1_3141_17358# vss nfet$261
Xnfet$254_5 m1_4005_21786# m1_4005_21786# vss vss m1_2843_21586# vss nfet$254
Xpfet$239_5 vdd m1_32817_25662# m1_32554_23922# m1_32330_25662# pfet$239
Xpfet$246_6 vdd m1_28470_16080# m1_28003_18030# m1_27031_17343# pfet$246
Xpfet$253_7 vdd vdd m1_n3541_23922# m1_n3184_24224# pfet$253
Xnfet$252_2 pd9 vss m1_26873_21786# vss nfet$252
Xnfet$245_1 m1_9015_17714# vss m1_6116_17343# vss nfet$245
Xpfet$251_4 vdd m1_n10452_25858# vdd m1_n4362_24346# pfet$251
Xpfet$228_108 vdd vdd m1_15454_18030# m1_15564_15778# pfet$228
Xnfet$247_13 m1_13198_17714# vss m1_16452_19550# vss nfet$247
Xpfet$230_9 vdd m1_9624_19404# m1_9624_19404# m1_9856_19850# m1_9418_19550# m1_9418_19550#
+ pfet$230
Xpfet$242_0 vdd vdd vdd m1_36073_22344# define define pfet$242
Xnfet$244_14 m1_17381_17714# m1_17381_17714# vss vss m1_21039_20470# vss nfet$244
Xnfet$269_11 m1_n10452_25858# vss m1_n4847_25662# vss nfet$269
Xpfet$227_97 vdd vdd m1_21590_21786# m1_24309_25858# pfet$227
Xpfet$227_86 vdd m1_28634_25662# m1_28371_23922# m1_28147_25662# pfet$227
Xpfet$227_75 vdd vdd m1_19644_25858# m1_14556_21786# pfet$227
Xpfet$227_64 vdd vdd m1_22522_24542# m1_20126_25858# pfet$227
Xpfet$227_53 vdd m1_20625_24224# m1_21729_25658# m1_19644_25858# pfet$227
Xpfet$227_42 vdd m1_11760_25858# vdd m1_13363_25658# pfet$227
Xnfet$249_8 m1_n7513_20152# vss m1_26676_16080# vss nfet$249
Xpfet$227_31 vdd m1_3273_23922# m1_3537_24542# m1_2912_25858# pfet$227
Xpfet$227_20 vdd vdd m1_4509_24346# m1_n7513_20152# pfet$227
Xnfet$268_0 m1_n3822_20130# m1_n3822_20130# m1_n4485_20152# m1_n4485_20152# m1_n3724_20470#
+ vss nfet$268
Xnfet$275_1 m1_n2543_20130# m1_n2543_20130# m1_n5227_20152# m1_n5227_20152# m1_n2445_20470#
+ vss nfet$275
Xnfet$241_26 m1_25912_25658# m1_25912_25658# vss vss m1_26371_25502# vss nfet$241
Xnfet$241_15 m1_25424_24346# m1_25424_24346# vss vss m1_24906_24542# vss nfet$241
Xnfet$247_5 m1_965_15478# vss m1_8137_20152# vss nfet$247
Xnfet$261_7 m1_5761_16080# m1_5761_16080# m1_5302_17714# m1_5302_17714# m1_5859_16398#
+ vss nfet$261
Xnfet$254_6 m1_4637_21786# m1_4637_21786# vss vss m1_3475_21586# vss nfet$254
Xpfet$239_6 vdd m1_34278_25658# m1_35071_24542# m1_32330_25662# pfet$239
Xpfet$246_7 vdd m1_27292_16202# m1_26807_17518# m1_27190_17836# pfet$246
Xpfet$253_8 vdd vdd m1_n2567_23922# m1_n7320_25516# pfet$253
.ends

.subckt pfet$295 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$293 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$314 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$312 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$296 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$294 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$313 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt nfet$311 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt asc_drive_buffer$3 vss in vdd out
Xpfet$295_0 vdd vdd m1_4002_n1060# m1_3466_n454# pfet$295
Xpfet$293_0 out out m1_4274_n1060# vdd m1_4274_n1060# out vdd vdd m1_4274_n1060# out
+ m1_4274_n1060# m1_4274_n1060# out m1_4274_n1060# vdd m1_4274_n1060# vdd m1_4274_n1060#
+ pfet$293
Xnfet$314_0 in vss m1_3466_n454# vss nfet$314
Xnfet$312_0 out out vss m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# m1_4274_n1060#
+ m1_4274_n1060# out m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# vss vss
+ nfet$312
Xpfet$296_0 vdd vdd m1_3466_n454# in pfet$296
Xpfet$294_0 m1_4274_n1060# vdd vdd m1_4274_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ vdd m1_4002_n1060# m1_4002_n1060# pfet$294
Xnfet$313_0 m1_3466_n454# vss m1_4002_n1060# vss nfet$313
Xnfet$311_0 m1_4274_n1060# vss m1_4002_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ m1_4274_n1060# vss m1_4002_n1060# vss nfet$311
.ends

.subckt asc_hysteresis_buffer$3 vss in vdd out
Xpfet$270_0 vdd vdd m1_884_42# m1_1156_42# pfet$270
Xnfet$287_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$287
Xnfet$285_0 m1_348_648# vss m1_884_42# vss nfet$285
Xpfet$268_0 vdd vdd m1_348_648# in pfet$268
Xpfet$266_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd
+ m1_884_42# m1_884_42# pfet$266
Xnfet$288_0 m1_1156_42# vss m1_884_42# vss nfet$288
Xnfet$286_0 in vss m1_348_648# vss nfet$286
Xnfet$284_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$284
Xpfet$269_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$269
Xpfet$267_0 vdd vdd m1_884_42# m1_348_648# pfet$267
.ends

.subckt xp_3_1_MUX$2 S0 S1 VDD VSS OUT_1 C_1 B_1 A_1
Xpfet$286_0 VDD A_1 m1_239_n318# m1_n432_458# pfet$286
Xpfet$286_2 VDD B_1 m1_239_n318# S0 pfet$286
Xpfet$286_1 VDD C_1 OUT_1 S1 pfet$286
Xpfet$286_3 VDD m1_239_n318# OUT_1 m1_n432_n1290# pfet$286
Xnfet$305_0 S1 VSS m1_n432_n1290# VSS nfet$305
Xnfet$305_1 S0 VSS m1_n432_458# VSS nfet$305
Xpfet$287_0 VDD VDD m1_n432_n1290# S1 pfet$287
Xpfet$287_1 VDD VDD m1_n432_458# S0 pfet$287
Xnfet$304_0 m1_n432_n1290# C_1 OUT_1 VSS nfet$304
Xnfet$304_1 m1_n432_458# B_1 m1_239_n318# VSS nfet$304
Xnfet$304_2 S1 m1_239_n318# OUT_1 VSS nfet$304
Xnfet$304_3 S0 A_1 m1_239_n318# VSS nfet$304
.ends

.subckt nfet$279 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$265 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.5u
.ends

.subckt nfet$280 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$262 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=4.55p ps=15.3u w=7u l=0.5u
.ends

.subckt pfet$261 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_954_0# w_n180_n88#
+ a_38_n60# a_n92_0# a_1058_n60# a_854_n60# a_342_0# a_138_0# a_650_n60#
X0 a_954_0# a_854_n60# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n60# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt nfet$278 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$260 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_954_0# w_n180_n88# a_854_n136#
+ a_n92_0# a_446_n136# a_650_n136# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt nfet$283 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$263 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$281 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pass1u05u$2 VDD VSS ind ins clkn clkp
Xpfet$263_0 VDD ind ins clkp pfet$263
Xnfet$281_0 clkn ind ins VSS nfet$281
.ends

.subckt pfet$264 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$282 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt inv1u05u$2 VDD in VSS out
Xpfet$264_0 VDD VDD out in pfet$264
Xnfet$282_0 in VSS out VSS nfet$282
.ends

.subckt xp_programmable_basic_pump$1 up vdd s1 s2 s3 s4 down out iref vss
Xnfet$279_8 down down vss vss m1_n8807_n11192# vss nfet$279
Xpfet$265_0 vdd s3 pass1u05u$2_5/ins vdd pfet$265
Xnfet$280_0 m1_n7879_n12170# pass1u05u$2_0/ins m1_n7879_n12170# out pass1u05u$2_0/ins
+ vss nfet$280
Xnfet$279_9 down down vss vss m1_n8807_n11192# vss nfet$279
Xpfet$265_1 vdd s2 pass1u05u$2_4/ins vdd pfet$265
Xnfet$280_1 m1_n7879_n12170# pass1u05u$2_0/ins m1_n7879_n12170# out pass1u05u$2_0/ins
+ vss nfet$280
Xpfet$262_20 vdd vdd vdd vdd pfet$262
Xpfet$265_2 vdd s1 pass1u05u$2_3/ins vdd pfet$265
Xnfet$280_2 vss down vss m1_n7879_n12170# down vss nfet$280
Xpfet$262_21 vdd vdd vdd vdd pfet$262
Xpfet$262_10 vdd vdd vdd vdd pfet$262
Xpfet$265_3 vdd s4 pass1u05u$2_7/ins vdd pfet$265
Xnfet$280_3 vss down vss m1_n7879_n12170# down vss nfet$280
Xpfet$262_22 vdd vdd vdd vdd pfet$262
Xpfet$262_11 vdd vdd vdd vdd pfet$262
Xnfet$280_4 vss down vss m1_n7879_n12170# down vss nfet$280
Xpfet$262_23 vdd vdd vdd vdd pfet$262
Xpfet$262_12 vdd vdd vdd vdd pfet$262
Xnfet$280_5 vss down vss m1_n7879_n12170# down vss nfet$280
Xpfet$262_13 vdd vdd vdd vdd pfet$262
Xnfet$280_6 m1_n7879_n12170# pass1u05u$2_0/ins m1_n7879_n12170# out pass1u05u$2_0/ins
+ vss nfet$280
Xpfet$261_0 vdd vdd m1_n4127_3649# vss vss m1_n4127_3649# vdd vss vdd vss vss vdd
+ m1_n4127_3649# vss pfet$261
Xpfet$262_14 vdd vdd vdd vdd pfet$262
Xnfet$280_7 m1_n7879_n12170# pass1u05u$2_0/ins m1_n7879_n12170# out pass1u05u$2_0/ins
+ vss nfet$280
Xpfet$262_15 vdd vdd vdd vdd pfet$262
Xpfet$261_1 m1_n5580_883# m1_n5580_883# out pass1u05u$2_5/ins pass1u05u$2_5/ins out
+ vdd pass1u05u$2_5/ins m1_n5580_883# pass1u05u$2_5/ins pass1u05u$2_5/ins m1_n5580_883#
+ out pass1u05u$2_5/ins pfet$261
Xnfet$280_8 vss vdd vss m1_n8144_n9165# vdd vss nfet$280
Xpfet$262_16 vdd vdd vdd vdd pfet$262
Xpfet$261_2 m1_n5580_883# m1_n5580_883# out pass1u05u$2_5/ins pass1u05u$2_5/ins out
+ vdd pass1u05u$2_5/ins m1_n5580_883# pass1u05u$2_5/ins pass1u05u$2_5/ins m1_n5580_883#
+ out pass1u05u$2_5/ins pfet$261
Xnfet$280_9 m1_n7216_n8262# iref m1_n7216_n8262# pass1u05u$2_7/ind iref vss nfet$280
Xpfet$262_17 vdd vdd vdd vdd pfet$262
Xpfet$261_3 m1_n5580_883# m1_n5580_883# out pass1u05u$2_5/ins pass1u05u$2_5/ins out
+ vdd pass1u05u$2_5/ins m1_n5580_883# pass1u05u$2_5/ins pass1u05u$2_5/ins m1_n5580_883#
+ out pass1u05u$2_5/ins pfet$261
Xnfet$280_10 m1_n8607_n8040# pass1u05u$2_1/ins m1_n8607_n8040# out pass1u05u$2_1/ins
+ vss nfet$280
Xnfet$278_10 pass1u05u$2_2/ins pass1u05u$2_2/ins m1_n7679_n8960# m1_n7679_n8960# out
+ vss nfet$278
Xpfet$262_18 vdd vdd vdd vdd pfet$262
Xpfet$261_4 m1_n5580_883# m1_n5580_883# out pass1u05u$2_5/ins pass1u05u$2_5/ins out
+ vdd pass1u05u$2_5/ins m1_n5580_883# pass1u05u$2_5/ins pass1u05u$2_5/ins m1_n5580_883#
+ out pass1u05u$2_5/ins pfet$261
Xnfet$280_11 m1_n8144_n9165# iref m1_n8144_n9165# iref iref vss nfet$280
Xnfet$278_0 pass1u05u$2_6/ins pass1u05u$2_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$278
Xpfet$261_5 m1_n4127_3649# m1_n4127_3649# pass1u05u$2_7/ind pass1u05u$2_7/ind pass1u05u$2_7/ind
+ pass1u05u$2_7/ind vdd pass1u05u$2_7/ind m1_n4127_3649# pass1u05u$2_7/ind pass1u05u$2_7/ind
+ m1_n4127_3649# pass1u05u$2_7/ind pass1u05u$2_7/ind pfet$261
Xnfet$278_11 vss vss vss vss vss vss nfet$278
Xnfet$280_12 vss down vss m1_n8607_n8040# down vss nfet$280
Xpfet$262_19 vdd vdd vdd vdd pfet$262
Xnfet$278_1 pass1u05u$2_6/ins pass1u05u$2_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$278
Xnfet$278_12 down down vss vss m1_n7679_n8960# vss nfet$278
Xnfet$280_13 vss vdd vss m1_n7216_n8262# vdd vss nfet$280
Xpfet$260_20 m1_n8156_628# m1_n8156_628# pass1u05u$2_7/ins out out vdd pass1u05u$2_7/ins
+ m1_n8156_628# pass1u05u$2_7/ins pass1u05u$2_7/ins m1_n8156_628# out pass1u05u$2_7/ins
+ pass1u05u$2_7/ins pfet$260
Xnfet$278_2 pass1u05u$2_6/ins pass1u05u$2_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$278
Xnfet$278_13 vss vss vss vss vss vss nfet$278
Xnfet$283_0 inv1u05u$2_2/out pass1u05u$2_1/ins vss vss nfet$283
Xnfet$280_14 m1_n8607_n8040# pass1u05u$2_1/ins m1_n8607_n8040# out pass1u05u$2_1/ins
+ vss nfet$280
Xpass1u05u$2_0 vdd vss iref pass1u05u$2_0/ins s3 inv1u05u$2_1/out pass1u05u$2
Xnfet$278_14 vss vss vss vss vss vss nfet$278
Xpfet$260_21 m1_n6703_2564# m1_n6703_2564# pass1u05u$2_4/ins out out vdd pass1u05u$2_4/ins
+ m1_n6703_2564# pass1u05u$2_4/ins pass1u05u$2_4/ins m1_n6703_2564# out pass1u05u$2_4/ins
+ pass1u05u$2_4/ins pfet$260
Xnfet$283_1 inv1u05u$2_3/out pass1u05u$2_2/ins vss vss nfet$283
Xnfet$278_3 vss vss vss vss vss vss nfet$278
Xpfet$260_10 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$260
Xpass1u05u$2_1 vdd vss iref pass1u05u$2_1/ins s2 inv1u05u$2_2/out pass1u05u$2
Xnfet$280_15 vss down vss m1_n8607_n8040# down vss nfet$280
Xpfet$260_22 m1_n8156_628# m1_n8156_628# pass1u05u$2_7/ins out out vdd pass1u05u$2_7/ins
+ m1_n8156_628# pass1u05u$2_7/ins pass1u05u$2_7/ins m1_n8156_628# out pass1u05u$2_7/ins
+ pass1u05u$2_7/ins pfet$260
Xnfet$278_4 pass1u05u$2_6/ins pass1u05u$2_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$278
Xpfet$260_11 vdd vdd up m1_n5450_4559# m1_n5450_4559# vdd up vdd up up vdd m1_n5450_4559#
+ up up pfet$260
Xnfet$278_15 vss vss vss vss vss vss nfet$278
Xnfet$283_2 inv1u05u$2_0/out pass1u05u$2_6/ins vss vss nfet$283
Xpass1u05u$2_2 vdd vss iref pass1u05u$2_2/ins s1 inv1u05u$2_3/out pass1u05u$2
Xpfet$260_23 m1_n8156_628# m1_n8156_628# pass1u05u$2_7/ins out out vdd pass1u05u$2_7/ins
+ m1_n8156_628# pass1u05u$2_7/ins pass1u05u$2_7/ins m1_n8156_628# out pass1u05u$2_7/ins
+ pass1u05u$2_7/ins pfet$260
Xnfet$283_3 inv1u05u$2_1/out pass1u05u$2_0/ins vss vss nfet$283
Xnfet$278_5 vss vss vss vss vss vss nfet$278
Xpfet$260_12 vdd vdd up m1_n6703_2564# m1_n6703_2564# vdd up vdd up up vdd m1_n6703_2564#
+ up up pfet$260
Xpass1u05u$2_3 vdd vss pass1u05u$2_7/ind pass1u05u$2_3/ins s1 inv1u05u$2_3/out pass1u05u$2
Xpfet$260_24 m1_n5450_4559# m1_n5450_4559# pass1u05u$2_3/ins out out vdd pass1u05u$2_3/ins
+ m1_n5450_4559# pass1u05u$2_3/ins pass1u05u$2_3/ins m1_n5450_4559# out pass1u05u$2_3/ins
+ pass1u05u$2_3/ins pfet$260
Xnfet$278_6 pass1u05u$2_6/ins pass1u05u$2_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$278
Xpfet$260_13 vdd vdd up m1_n6703_2564# m1_n6703_2564# vdd up vdd up up vdd m1_n6703_2564#
+ up up pfet$260
Xinv1u05u$2_0 vdd s4 vss inv1u05u$2_0/out inv1u05u$2
Xpass1u05u$2_4 vdd vss pass1u05u$2_7/ind pass1u05u$2_4/ins s2 inv1u05u$2_2/out pass1u05u$2
Xpfet$260_25 m1_n6703_2564# m1_n6703_2564# pass1u05u$2_4/ins out out vdd pass1u05u$2_4/ins
+ m1_n6703_2564# pass1u05u$2_4/ins pass1u05u$2_4/ins m1_n6703_2564# out pass1u05u$2_4/ins
+ pass1u05u$2_4/ins pfet$260
Xinv1u05u$2_1 vdd s3 vss inv1u05u$2_1/out inv1u05u$2
Xnfet$278_7 pass1u05u$2_6/ins pass1u05u$2_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$278
Xpfet$260_14 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$260
Xpass1u05u$2_5 vdd vss pass1u05u$2_7/ind pass1u05u$2_5/ins s3 inv1u05u$2_1/out pass1u05u$2
Xnfet$278_8 pass1u05u$2_6/ins pass1u05u$2_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$278
Xpfet$260_15 m1_n8156_628# m1_n8156_628# pass1u05u$2_7/ins out out vdd pass1u05u$2_7/ins
+ m1_n8156_628# pass1u05u$2_7/ins pass1u05u$2_7/ins m1_n8156_628# out pass1u05u$2_7/ins
+ pass1u05u$2_7/ins pfet$260
Xinv1u05u$2_2 vdd s2 vss inv1u05u$2_2/out inv1u05u$2
Xpass1u05u$2_6 vdd vss iref pass1u05u$2_6/ins s4 inv1u05u$2_0/out pass1u05u$2
Xinv1u05u$2_3 vdd s1 vss inv1u05u$2_3/out inv1u05u$2
Xnfet$278_9 pass1u05u$2_6/ins pass1u05u$2_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$278
Xpfet$260_16 m1_n8156_628# m1_n8156_628# pass1u05u$2_7/ins out out vdd pass1u05u$2_7/ins
+ m1_n8156_628# pass1u05u$2_7/ins pass1u05u$2_7/ins m1_n8156_628# out pass1u05u$2_7/ins
+ pass1u05u$2_7/ins pfet$260
Xpass1u05u$2_7 vdd vss pass1u05u$2_7/ind pass1u05u$2_7/ins s4 inv1u05u$2_0/out pass1u05u$2
Xpfet$260_17 m1_n8156_628# m1_n8156_628# pass1u05u$2_7/ins out out vdd pass1u05u$2_7/ins
+ m1_n8156_628# pass1u05u$2_7/ins pass1u05u$2_7/ins m1_n8156_628# out pass1u05u$2_7/ins
+ pass1u05u$2_7/ins pfet$260
Xpfet$260_18 m1_n8156_628# m1_n8156_628# pass1u05u$2_7/ins out out vdd pass1u05u$2_7/ins
+ m1_n8156_628# pass1u05u$2_7/ins pass1u05u$2_7/ins m1_n8156_628# out pass1u05u$2_7/ins
+ pass1u05u$2_7/ins pfet$260
Xnfet$279_10 vss vss vss vss vss vss nfet$279
Xpfet$262_0 vdd vdd vdd vdd pfet$262
Xpfet$260_19 m1_n8156_628# m1_n8156_628# pass1u05u$2_7/ins out out vdd pass1u05u$2_7/ins
+ m1_n8156_628# pass1u05u$2_7/ins pass1u05u$2_7/ins m1_n8156_628# out pass1u05u$2_7/ins
+ pass1u05u$2_7/ins pfet$260
Xnfet$279_11 vss vss vss vss vss vss nfet$279
Xpfet$262_1 vdd vdd vdd vdd pfet$262
Xnfet$279_12 vss vss vss vss vss vss nfet$279
Xpfet$262_2 vdd vdd vdd vdd pfet$262
Xnfet$279_13 vss vss vss vss vss vss nfet$279
Xpfet$262_3 vdd vdd vdd vdd pfet$262
Xpfet$260_0 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$260
Xpfet$262_4 vdd vdd vdd vdd pfet$262
Xpfet$260_1 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$260
Xnfet$279_0 down down vss vss m1_n8807_n11192# vss nfet$279
Xpfet$260_2 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$260
Xpfet$262_5 vdd vdd vdd vdd pfet$262
Xnfet$279_1 down down vss vss m1_n8807_n11192# vss nfet$279
Xpfet$262_6 vdd vdd vdd vdd pfet$262
Xpfet$260_3 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$260
Xnfet$279_2 down down vss vss m1_n8807_n11192# vss nfet$279
Xpfet$260_4 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$260
Xpfet$262_7 vdd vdd vdd vdd pfet$262
Xnfet$279_3 down down vss vss m1_n8807_n11192# vss nfet$279
Xpfet$262_8 vdd vdd vdd vdd pfet$262
Xpfet$260_5 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$260
Xnfet$279_4 vss vss vss vss vss vss nfet$279
Xpfet$260_6 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$260
Xpfet$262_9 vdd vdd vdd vdd pfet$262
Xnfet$279_5 vss vss vss vss vss vss nfet$279
Xpfet$260_7 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$260
Xnfet$279_6 down down vss vss m1_n8807_n11192# vss nfet$279
Xpfet$260_8 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$260
Xnfet$279_7 down down vss vss m1_n8807_n11192# vss nfet$279
Xpfet$260_9 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$260
.ends

.subckt asc_dual_psd_def_20250809$2 vdd vss pd1 pd2 pd3 pd4 pd5 pd6 pd7 pd8 pd9 fout
+ sd1 sd2 sd3 sd4 sd5 sd6 sd7 sd8 sd9 fin define
Xnfet$242_80 m1_28147_25662# m1_28991_24224# m1_30095_25658# vss nfet$242
Xnfet$245_2 m1_6275_17836# m1_7555_16080# m1_7088_18030# vss nfet$245
Xpfet$251_5 vdd vdd m1_n10308_24542# m1_n9952_24224# pfet$251
Xpfet$228_109 vdd vdd m1_10299_17343# m1_13198_17714# pfet$228
Xnfet$247_14 m1_21564_17714# vss m1_23486_19550# vss nfet$247
Xnfet$250_0 m1_n10452_25858# vss m1_n1271_25858# vss nfet$250
Xpfet$242_1 vdd m1_35837_22102# m1_35837_22102# m1_36073_22344# fout fout pfet$242
Xpfet$235_0 vdd vdd m1_n647_25662# m1_n789_25858# pfet$235
Xnfet$244_15 m1_21564_17714# m1_21564_17714# vss vss m1_24556_20470# vss nfet$244
Xnfet$269_12 m1_n10452_25858# vss m1_n5571_25662# vss nfet$269
Xpfet$232_10 vdd vdd m1_27031_17343# m1_n10452_25858# pfet$232
Xpfet$227_65 vdd vdd m1_18073_21786# m1_20126_25858# pfet$227
Xpfet$227_54 vdd vdd m1_24808_24224# m1_24188_23922# pfet$227
Xpfet$227_43 vdd vdd m1_12805_21786# pd5 pfet$227
Xnfet$245_80 m1_18824_17836# m1_19747_15778# m1_18926_16202# vss nfet$245
Xnfet$249_9 m1_n10452_25858# vss m1_27031_17343# vss nfet$249
Xpfet$227_32 vdd vdd m1_7720_24542# m1_8076_24224# pfet$227
Xpfet$227_21 vdd m1_7456_23922# m1_7720_24542# m1_7095_25858# pfet$227
Xpfet$227_10 vdd m1_8076_24224# m1_9180_25658# m1_7095_25858# pfet$227
Xnfet$268_1 m1_n1927_20274# m1_n1927_20274# vss vss m1_n2445_20470# vss nfet$268
Xnfet$241_27 m1_12875_24346# m1_12875_24346# vss vss m1_12357_24542# vss nfet$241
Xpfet$227_98 vdd m1_30095_25658# m1_30888_24542# m1_28147_25662# pfet$227
Xpfet$227_87 vdd vdd m1_28147_25662# m1_28010_25858# pfet$227
Xpfet$227_76 vdd m1_20005_23922# m1_20269_24542# m1_19644_25858# pfet$227
Xnfet$241_16 m1_24808_24224# m1_24808_24224# m1_24452_24542# m1_24452_24542# m1_24906_24542#
+ vss nfet$241
Xnfet$254_7 m1_488_21786# m1_488_21786# vss vss m1_n674_21586# vss nfet$254
Xnfet$247_6 m1_9015_17714# vss m1_12935_19550# vss nfet$247
Xnfet$261_8 m1_3015_15778# m1_3015_15778# m1_2905_18030# m1_2905_18030# m1_3141_17358#
+ vss nfet$261
Xpfet$239_7 vdd m1_32554_23922# m1_32818_24542# m1_32193_25858# pfet$239
Xpfet$253_9 vdd vdd m1_n4464_25980# m1_n4623_25487# pfet$253
Xnfet$242_81 m1_n7513_20152# vss m1_25424_24346# vss nfet$242
Xnfet$242_70 m1_21590_21786# vss m1_28010_25858# vss nfet$242
Xnfet$245_3 m1_n7513_20152# vss m1_9944_16080# vss nfet$245
Xnfet$247_15 m1_17697_15478# vss m1_22205_20152# vss nfet$247
Xpfet$251_6 vdd m1_n10308_24542# vdd m1_n9336_24346# pfet$251
Xpfet$227_110 vdd m1_11903_24542# vdd m1_12875_24346# pfet$227
Xpfet$235_10 vdd vdd m1_35071_24542# m1_32675_25947# pfet$235
Xnfet$243_0 m1_n1133_21590# m1_n1133_21590# m1_354_22513# m1_354_22513# m1_n674_21586#
+ vss nfet$243
Xpfet$235_1 vdd vdd m1_n1134_25662# m1_n1271_25858# pfet$235
Xnfet$250_1 m1_n789_25858# vss m1_n647_25662# vss nfet$250
Xpfet$228_0 vdd vdd m1_12355_15778# m1_9485_17714# pfet$228
Xnfet$244_16 m1_23486_19550# m1_23486_19550# vss vss m1_23924_20470# vss nfet$244
Xnfet$269_13 fin vss m1_n4623_25487# vss nfet$269
Xpfet$232_11 vdd vdd m1_26807_17518# m1_26217_17714# pfet$232
Xnfet$245_81 m1_13198_17714# vss m1_10299_17343# vss nfet$245
Xnfet$245_70 m1_n7513_20152# vss m1_18310_16080# vss nfet$245
Xpfet$227_99 vdd vdd m1_26705_24542# m1_24309_25858# pfet$227
Xpfet$227_88 vdd vdd m1_28634_25662# m1_28492_25858# pfet$227
Xpfet$227_77 vdd vdd m1_20269_24542# m1_20625_24224# pfet$227
Xpfet$227_66 vdd vdd m1_15461_25858# m1_11039_21786# pfet$227
Xpfet$227_55 vdd m1_24451_25662# m1_24188_23922# m1_23964_25662# pfet$227
Xnfet$241_17 m1_20625_24224# m1_20625_24224# m1_20269_24542# m1_20269_24542# m1_20723_24542#
+ vss nfet$241
Xpfet$227_44 vdd m1_15943_25858# vdd m1_17546_25658# pfet$227
Xpfet$227_33 vdd vdd m1_7522_21786# m1_7577_25858# pfet$227
Xpfet$227_22 vdd vdd m1_3537_24542# m1_3893_24224# pfet$227
Xpfet$227_11 vdd vdd m1_7719_25662# m1_7577_25858# pfet$227
Xnfet$268_2 m1_n3206_20274# m1_n3206_20274# vss vss m1_n3724_20470# vss nfet$268
Xnfet$261_9 m1_2194_16202# m1_2194_16202# vss vss m1_1676_16398# vss nfet$261
Xnfet$254_8 m1_25739_21786# m1_25739_21786# vss vss m1_24577_21586# vss nfet$254
Xnfet$247_7 m1_5148_15478# vss m1_11654_20152# vss nfet$247
Xnfet$273_0 m1_n8283_20611# vss m1_n8283_19850# vss nfet$273
Xpfet$258_0 vdd vdd vdd m1_n5019_19550# m1_n4485_20152# m1_n4485_20152# pfet$258
Xnfet$242_82 m1_11415_25662# m1_12259_24224# m1_13363_25658# vss nfet$242
Xnfet$242_71 m1_28147_25662# m1_28371_23922# m1_28635_24542# vss nfet$242
Xnfet$242_60 pd6 vss m1_16322_21786# vss nfet$242
Xnfet$245_4 m1_10299_17343# m1_10560_16202# m1_10075_17518# vss nfet$245
Xnfet$247_16 m1_17381_17714# vss m1_19969_19550# vss nfet$247
Xpfet$251_7 vdd vdd m1_n10452_25858# m1_n4978_24224# pfet$251
Xpfet$235_11 vdd vdd m1_32817_25662# m1_32675_25947# pfet$235
Xpfet$227_100 vdd vdd m1_29607_24346# m1_n7513_20152# pfet$227
Xnfet$243_1 m1_n1263_21786# m1_n1263_21786# m1_354_22513# m1_354_22513# m1_n42_21586#
+ vss nfet$243
Xnfet$250_2 m1_n1271_25858# vss m1_n1134_25662# vss nfet$250
Xpfet$228_1 vdd vdd m1_11381_15778# m1_11738_16080# pfet$228
Xpfet$235_2 vdd vdd m1_n1271_25858# m1_n10452_25858# pfet$235
Xnfet$244_17 m1_12935_19550# m1_12935_19550# vss vss m1_13373_20470# vss nfet$244
Xpfet$240_0 vdd vdd m1_n1263_21786# pd1 pfet$240
Xpfet$232_12 vdd vdd m1_26676_16080# m1_n7513_20152# pfet$232
Xnfet$245_82 m1_10299_17343# vss m1_10458_17836# vss nfet$245
Xnfet$245_71 m1_14641_17836# m1_15921_16080# m1_15454_18030# vss nfet$245
Xnfet$245_60 m1_18665_17343# vss m1_18824_17836# vss nfet$245
Xpfet$227_89 vdd vdd m1_19839_21786# pd7 pfet$227
Xpfet$227_78 vdd m1_20269_24542# vdd m1_21241_24346# pfet$227
Xpfet$227_67 vdd m1_15822_23922# m1_16086_24542# m1_15461_25858# pfet$227
Xpfet$227_56 vdd m1_24808_24224# m1_25912_25658# m1_23827_25858# pfet$227
Xpfet$227_45 vdd vdd m1_16442_24224# m1_15822_23922# pfet$227
Xpfet$227_34 vdd m1_9180_25658# m1_9973_24542# m1_7232_25662# pfet$227
Xpfet$227_23 vdd m1_3537_24542# vdd m1_4509_24346# pfet$227
Xpfet$227_12 vdd m1_7577_25858# vdd m1_9180_25658# pfet$227
Xnfet$268_3 m1_n6973_21481# m1_n6973_21481# m1_n6839_20152# m1_n6839_20152# m1_n6282_20470#
+ vss nfet$268
Xnfet$241_18 m1_21241_24346# m1_21241_24346# vss vss m1_20723_24542# vss nfet$241
Xnfet$254_9 m1_25107_21786# m1_25107_21786# vss vss m1_23945_21586# vss nfet$254
Xnfet$273_1 m1_n7513_20152# m1_n8283_19850# vss vss nfet$273
Xnfet$247_8 m1_n7383_17599# vss m1_n1133_19550# vss nfet$247
Xnfet$266_0 m1_n10452_25858# m1_n10452_25858# m1_n7186_25858# m1_n7186_25858# m1_n6629_25502#
+ vss nfet$266
Xnfet$242_72 m1_23827_25858# m1_25912_25658# m1_26705_24542# vss nfet$242
Xnfet$242_61 m1_23964_25662# m1_24808_24224# m1_25912_25658# vss nfet$242
Xnfet$242_50 m1_n7513_20152# vss m1_21241_24346# vss nfet$242
Xnfet$245_5 m1_10458_17836# m1_11738_16080# m1_11271_18030# vss nfet$245
Xnfet$247_17 m1_21880_15478# vss m1_25722_20152# vss nfet$247
Xpfet$235_12 vdd vdd m1_32193_25858# m1_25107_21786# pfet$235
Xpfet$227_101 vdd vdd m1_28010_25858# m1_21590_21786# pfet$227
Xnfet$243_2 m1_9288_21786# m1_9288_21786# m1_9645_21447# m1_9645_21447# m1_10509_21586#
+ vss nfet$243
Xnfet$250_3 m1_n7513_20152# vss m1_326_24346# vss nfet$250
Xpfet$235_3 vdd vdd m1_1607_24542# m1_n789_25858# pfet$235
Xpfet$228_2 vdd m1_12355_15778# m1_11738_16080# m1_10458_17836# pfet$228
Xpfet$240_1 vdd vdd m1_2254_21786# pd2 pfet$240
Xpfet$233_0 vdd vdd m1_2384_19550# m1_n3534_17714# pfet$233
Xpfet$232_13 vdd vdd m1_25747_17714# m1_26217_17714# pfet$232
Xpfet$227_79 vdd m1_17546_25658# m1_18339_24542# m1_15598_25662# pfet$227
Xpfet$227_68 vdd vdd m1_16086_24542# m1_16442_24224# pfet$227
Xpfet$227_57 vdd vdd m1_24451_25662# m1_24309_25858# pfet$227
Xpfet$227_46 vdd m1_16442_24224# m1_17546_25658# m1_15461_25858# pfet$227
Xnfet$245_72 m1_17851_17714# vss m1_18441_17518# vss nfet$245
Xnfet$245_61 m1_20104_16080# vss m1_19747_15778# vss nfet$245
Xnfet$245_50 m1_25747_17714# vss m1_22848_17343# vss nfet$245
Xpfet$227_35 vdd m1_7720_24542# vdd m1_8692_24346# pfet$227
Xpfet$227_24 vdd vdd m1_5790_24542# m1_3394_25858# pfet$227
Xpfet$227_13 vdd vdd m1_12259_24224# m1_11639_23922# pfet$227
Xnfet$268_4 m1_2590_19404# m1_2590_19404# vss vss m1_n2445_21430# vss nfet$268
Xnfet$241_19 m1_21729_25658# m1_21729_25658# vss vss m1_22188_25502# vss nfet$241
Xnfet$247_9 m1_25747_17714# vss m1_27003_19550# vss nfet$247
Xnfet$259_0 m1_34093_22102# vss fout vss nfet$259
Xnfet$273_2 m1_n8145_21908# vss m1_n8283_20611# vss nfet$273
Xnfet$266_1 m1_n6111_25858# m1_n6111_25858# vss vss m1_n6629_25502# vss nfet$266
Xnfet$242_73 m1_24309_25858# vss m1_21590_21786# vss nfet$242
Xnfet$242_62 m1_24188_23922# vss m1_24808_24224# vss nfet$242
Xnfet$242_51 m1_19644_25858# m1_21729_25658# m1_22522_24542# vss nfet$242
Xnfet$242_40 m1_15598_25662# m1_16442_24224# m1_17546_25658# vss nfet$242
Xnfet$245_6 m1_6116_17343# vss m1_6275_17836# vss nfet$245
Xpfet$235_13 vdd vdd m1_33790_24346# m1_n7513_20152# pfet$235
Xpfet$227_102 vdd m1_28371_23922# m1_28635_24542# m1_28010_25858# pfet$227
Xnfet$243_3 m1_9418_21590# m1_9418_21590# m1_9645_21447# m1_9645_21447# m1_9877_21586#
+ vss nfet$243
Xnfet$250_4 m1_n789_25858# vss m1_1607_24542# vss nfet$250
Xpfet$235_4 vdd vdd m1_488_21786# m1_n789_25858# pfet$235
Xpfet$228_3 vdd m1_11381_15778# m1_10560_16202# m1_10299_17343# pfet$228
Xnfet$241_0 m1_4509_24346# m1_4509_24346# vss vss m1_3991_24542# vss nfet$241
Xpfet$240_2 vdd vdd m1_26873_21786# pd9 pfet$240
Xpfet$233_1 vdd vdd m1_4620_20152# m1_n3218_15478# pfet$233
Xpfet$227_69 vdd vdd m1_12875_24346# m1_n7513_20152# pfet$227
Xpfet$227_58 vdd vdd m1_23964_25662# m1_23827_25858# pfet$227
Xpfet$227_47 vdd vdd m1_15943_25858# m1_17058_24346# pfet$227
Xnfet$245_73 m1_13668_17714# vss m1_16538_15778# vss nfet$245
Xnfet$245_62 m1_18665_17343# m1_20721_15778# m1_20104_16080# vss nfet$245
Xnfet$245_51 m1_n7513_20152# vss m1_22493_16080# vss nfet$245
Xpfet$227_36 vdd vdd m1_8692_24346# m1_n7513_20152# pfet$227
Xpfet$227_25 vdd vdd m1_4005_21786# m1_3394_25858# pfet$227
Xpfet$227_14 vdd vdd m1_11902_25662# m1_11760_25858# pfet$227
Xnfet$245_40 m1_n2250_17343# m1_n194_15778# m1_n811_16080# vss nfet$245
Xnfet$268_5 m1_6107_19404# m1_6107_19404# m1_n5227_21418# m1_n5227_21418# m1_n2445_21430#
+ vss nfet$268
Xnfet$273_3 m1_n8283_19850# m1_n8283_20611# vss vss nfet$273
Xnfet$242_63 m1_14556_21786# vss m1_19644_25858# vss nfet$242
Xnfet$242_52 m1_20126_25858# vss m1_22522_24542# vss nfet$242
Xnfet$242_41 pd5 vss m1_12805_21786# vss nfet$242
Xnfet$242_30 m1_n7513_20152# vss m1_17058_24346# vss nfet$242
Xpfet$228_90 vdd m1_19747_15778# m1_18926_16202# m1_18665_17343# pfet$228
Xnfet$242_74 pd8 vss m1_23356_21786# vss nfet$242
Xnfet$245_7 m1_9485_17714# vss m1_10075_17518# vss nfet$245
Xpfet$256_0 vdd m1_n6380_21786# m1_n6380_21786# m1_n5019_19550# m1_n5227_20152# m1_n5227_20152#
+ pfet$256
Xnfet$271_0 m1_n10933_25858# m1_n8848_25658# m1_n8055_24542# vss nfet$271
Xpfet$227_103 vdd vdd m1_28635_24542# m1_28991_24224# pfet$227
Xnfet$250_5 m1_n789_25858# vss m1_488_21786# vss nfet$250
Xpfet$235_5 vdd vdd m1_326_24346# m1_n7513_20152# pfet$235
Xpfet$228_4 vdd m1_9485_17714# vdd m1_10560_16202# pfet$228
Xnfet$243_4 m1_5901_21590# m1_5901_21590# m1_7388_22513# m1_7388_22513# m1_6360_21586#
+ vss nfet$243
Xnfet$241_1 m1_3893_24224# m1_3893_24224# m1_3537_24542# m1_3537_24542# m1_3991_24542#
+ vss nfet$241
Xpfet$233_2 vdd vdd m1_1103_20152# m1_n7401_15478# pfet$233
Xpfet$227_59 vdd vdd m1_16322_21786# pd6 pfet$227
Xpfet$227_48 vdd m1_16085_25662# m1_15822_23922# m1_15598_25662# pfet$227
Xnfet$245_74 m1_14482_17343# vss m1_14641_17836# vss nfet$245
Xnfet$245_63 m1_13668_17714# vss m1_14258_17518# vss nfet$245
Xnfet$245_52 m1_23007_17836# m1_24287_16080# m1_23820_18030# vss nfet$245
Xpfet$227_37 vdd vdd m1_9973_24542# m1_7577_25858# pfet$227
Xpfet$227_26 vdd m1_4997_25658# m1_5790_24542# m1_3049_25662# pfet$227
Xpfet$227_15 vdd m1_11902_25662# m1_11639_23922# m1_11415_25662# pfet$227
Xnfet$245_30 sd6 vss m1_5148_15478# vss nfet$245
Xnfet$245_41 m1_n2091_17836# m1_n1168_15778# m1_n1989_16202# vss nfet$245
Xnfet$268_6 m1_n5764_21786# m1_n5764_21786# vss vss m1_n6282_21430# vss nfet$268
Xpfet$228_91 vdd m1_24287_16080# m1_23820_18030# m1_22848_17343# pfet$228
Xpfet$228_80 vdd vdd m1_15564_15778# m1_15921_16080# pfet$228
Xnfet$242_75 m1_28371_23922# vss m1_28991_24224# vss nfet$242
Xnfet$242_64 m1_19644_25858# vss m1_19781_25662# vss nfet$242
Xnfet$242_53 m1_23827_25858# m1_24451_25662# m1_24188_23922# vss nfet$242
Xnfet$242_42 m1_15943_25858# vss m1_16085_25662# vss nfet$242
Xnfet$242_31 m1_15943_25858# vss m1_18339_24542# vss nfet$242
Xnfet$242_20 pd3 vss m1_5771_21786# vss nfet$242
Xnfet$245_8 m1_7555_16080# vss m1_7198_15778# vss nfet$245
Xnfet$264_0 m1_n6274_17836# m1_n4994_16080# m1_n5461_18030# vss nfet$264
Xnfet$271_1 m1_n10796_25662# m1_n10572_23922# m1_n10308_24542# vss nfet$271
Xpfet$256_1 vdd vdd vdd m1_n5019_22344# m1_n4485_21904# m1_n4485_21904# pfet$256
Xpfet$249_0 vdd m1_n10309_25662# m1_n10572_23922# m1_n10796_25662# pfet$249
Xpfet$227_104 vdd m1_25912_25658# m1_26705_24542# m1_23964_25662# pfet$227
Xnfet$250_6 m1_n910_23922# vss m1_n290_24224# vss nfet$250
Xpfet$235_6 vdd vdd m1_n290_24224# m1_n910_23922# pfet$235
Xnfet$243_5 m1_2254_21786# m1_2254_21786# m1_3871_22513# m1_3871_22513# m1_3475_21586#
+ vss nfet$243
Xpfet$228_5 vdd m1_7198_15778# m1_6377_16202# m1_6116_17343# pfet$228
Xnfet$241_2 m1_4997_25658# m1_4997_25658# vss vss m1_5456_25502# vss nfet$241
Xpfet$233_3 vdd vdd m1_5901_19550# m1_649_17714# pfet$233
Xnfet$245_75 sd3 vss m1_17697_15478# vss nfet$245
Xnfet$245_64 m1_13668_17714# vss m1_13198_17714# vss nfet$245
Xnfet$245_53 m1_22848_17343# vss m1_23007_17836# vss nfet$245
Xnfet$245_31 m1_1933_17343# m1_3989_15778# m1_3372_16080# vss nfet$245
Xnfet$245_20 m1_1119_17714# vss m1_1709_17518# vss nfet$245
Xnfet$245_42 m1_n811_16080# vss m1_n1168_15778# vss nfet$245
Xpfet$231_0 vdd vdd m1_n1133_21590# m1_n1263_21786# pfet$231
Xpfet$227_49 vdd m1_20126_25858# vdd m1_21729_25658# pfet$227
Xpfet$227_38 vdd vdd m1_16085_25662# m1_15943_25858# pfet$227
Xpfet$227_27 vdd vdd m1_11278_25858# m1_7522_21786# pfet$227
Xpfet$227_16 vdd vdd m1_5771_21786# pd3 pfet$227
Xnfet$268_7 m1_n3822_21786# m1_n3822_21786# m1_n4485_21904# m1_n4485_21904# m1_n3724_21430#
+ vss nfet$268
Xpfet$228_92 vdd m1_15454_18030# vdd m1_14127_16080# pfet$228
Xpfet$228_81 vdd vdd m1_13668_17714# m1_14127_16080# pfet$228
Xpfet$228_70 vdd vdd m1_18824_17836# m1_18665_17343# pfet$228
Xnfet$242_76 m1_28492_25858# vss m1_28634_25662# vss nfet$242
Xnfet$242_65 m1_28492_25858# vss m1_25107_21786# vss nfet$242
Xnfet$242_54 m1_24309_25858# vss m1_24451_25662# vss nfet$242
Xnfet$242_43 m1_15461_25858# vss m1_15598_25662# vss nfet$242
Xnfet$242_32 m1_15461_25858# m1_17546_25658# m1_18339_24542# vss nfet$242
Xnfet$242_21 m1_11278_25858# m1_11902_25662# m1_11639_23922# vss nfet$242
Xnfet$242_10 m1_7577_25858# vss m1_9973_24542# vss nfet$242
Xnfet$245_9 sd5 vss m1_9331_15478# vss nfet$245
Xnfet$257_0 m1_31535_22102# m1_32818_21586# vss vss nfet$257
Xnfet$264_1 m1_n6433_17343# m1_n4377_15778# m1_n4994_16080# vss nfet$264
Xnfet$271_2 m1_n10933_25858# m1_n10309_25662# m1_n10572_23922# vss nfet$271
Xpfet$256_2 vdd m1_n5764_21786# m1_n5764_21786# m1_n5019_22344# m1_n5227_21418# m1_n5227_21418#
+ pfet$256
Xpfet$249_1 vdd m1_n9952_24224# m1_n8848_25658# m1_n10933_25858# pfet$249
Xpfet$227_105 vdd vdd m1_30888_24542# m1_28492_25858# pfet$227
Xnfet$250_7 m1_25107_21786# vss m1_32193_25858# vss nfet$250
Xnfet$243_6 m1_2384_21590# m1_2384_21590# m1_3871_22513# m1_3871_22513# m1_2843_21586#
+ vss nfet$243
Xpfet$235_7 vdd vdd m1_32330_25662# m1_32193_25858# pfet$235
Xpfet$228_6 vdd vdd m1_7198_15778# m1_7555_16080# pfet$228
Xnfet$241_3 m1_4509_24346# m1_4509_24346# m1_3394_25858# m1_3394_25858# m1_5456_25502#
+ vss nfet$241
Xpfet$233_4 vdd vdd m1_12935_19550# m1_9015_17714# pfet$233
Xnfet$250_10 m1_32675_25947# vss m1_35071_24542# vss nfet$250
Xnfet$245_76 m1_14482_17343# m1_16538_15778# m1_15921_16080# vss nfet$245
Xnfet$245_65 m1_14482_17343# m1_14743_16202# m1_14258_17518# vss nfet$245
Xnfet$245_54 m1_22848_17343# m1_23109_16202# m1_22624_17518# vss nfet$245
Xnfet$245_32 m1_2092_17836# m1_3015_15778# m1_2194_16202# vss nfet$245
Xnfet$245_21 m1_1933_17343# m1_2194_16202# m1_1709_17518# vss nfet$245
Xnfet$245_10 m1_11738_16080# vss m1_11381_15778# vss nfet$245
Xnfet$245_43 sd8 vss m1_n3218_15478# vss nfet$245
Xpfet$231_1 vdd vdd m1_11671_21786# m1_11039_21786# pfet$231
Xpfet$227_39 vdd vdd m1_15598_25662# m1_15461_25858# pfet$227
Xnfet$261_20 m1_22493_16080# m1_22493_16080# m1_22034_17714# m1_22034_17714# m1_22591_16398#
+ vss nfet$261
Xpfet$227_28 vdd m1_11639_23922# m1_11903_24542# m1_11278_25858# pfet$227
Xpfet$227_17 vdd vdd m1_7577_25858# m1_8692_24346# pfet$227
Xnfet$268_8 m1_9624_19404# m1_9624_19404# vss vss m1_n3724_21430# vss nfet$268
Xpfet$228_93 vdd m1_23820_18030# vdd m1_22493_16080# pfet$228
Xpfet$228_82 vdd m1_13668_17714# vdd m1_14743_16202# pfet$228
Xpfet$228_71 vdd vdd m1_19747_15778# m1_20104_16080# pfet$228
Xpfet$228_60 vdd vdd m1_n194_15778# m1_n3064_17714# pfet$228
Xnfet$242_77 m1_28010_25858# vss m1_28147_25662# vss nfet$242
Xnfet$242_66 m1_28010_25858# m1_30095_25658# m1_30888_24542# vss nfet$242
Xnfet$242_55 m1_23827_25858# vss m1_23964_25662# vss nfet$242
Xnfet$242_44 m1_15822_23922# vss m1_16442_24224# vss nfet$242
Xnfet$242_33 m1_11760_25858# vss m1_14156_24542# vss nfet$242
Xnfet$242_22 m1_11760_25858# vss m1_11902_25662# vss nfet$242
Xnfet$242_11 m1_7522_21786# vss m1_11278_25858# vss nfet$242
Xnfet$264_2 m1_n6274_17836# m1_n5351_15778# m1_n6172_16202# vss nfet$264
Xnfet$271_3 m1_n10796_25662# m1_n9952_24224# m1_n8848_25658# vss nfet$271
Xpfet$249_2 vdd m1_n4362_24346# m1_n4847_25662# m1_n4464_25980# pfet$249
Xpfet$227_106 vdd vdd m1_25107_21786# m1_28492_25858# pfet$227
Xnfet$250_8 m1_32193_25858# vss m1_32330_25662# vss nfet$250
Xnfet$243_7 m1_5771_21786# m1_5771_21786# m1_7388_22513# m1_7388_22513# m1_6992_21586#
+ vss nfet$243
Xpfet$235_8 vdd vdd m1_33174_24224# m1_32554_23922# pfet$235
Xpfet$228_7 vdd vdd m1_6275_17836# m1_6116_17343# pfet$228
Xpfet$254_0 vdd vdd m1_n7186_25858# m1_n10452_25858# pfet$254
Xnfet$241_4 m1_12259_24224# m1_12259_24224# m1_11903_24542# m1_11903_24542# m1_12357_24542#
+ vss nfet$241
Xpfet$233_5 vdd vdd m1_8137_20152# m1_965_15478# pfet$233
Xnfet$250_11 m1_32554_23922# vss m1_33174_24224# vss nfet$250
Xpfet$231_2 vdd vdd m1_12935_21590# m1_12805_21786# pfet$231
Xnfet$245_77 sd4 vss m1_13514_15478# vss nfet$245
Xnfet$245_66 m1_n7513_20152# vss m1_14127_16080# vss nfet$245
Xnfet$261_21 m1_14127_16080# m1_14127_16080# vss vss m1_15690_17358# vss nfet$261
Xnfet$245_55 m1_22034_17714# vss m1_24904_15778# vss nfet$245
Xnfet$245_44 m1_n2091_17836# m1_n811_16080# m1_n1278_18030# vss nfet$245
Xpfet$227_29 vdd vdd m1_11903_24542# m1_12259_24224# pfet$227
Xpfet$227_18 vdd vdd m1_11415_25662# m1_11278_25858# pfet$227
Xnfet$245_33 sd7 vss m1_965_15478# vss nfet$245
Xnfet$261_10 m1_1578_16080# m1_1578_16080# m1_1119_17714# m1_1119_17714# m1_1676_16398#
+ vss nfet$261
Xnfet$245_22 m1_6116_17343# m1_6377_16202# m1_5892_17518# vss nfet$245
Xnfet$245_11 m1_10299_17343# m1_12355_15778# m1_11738_16080# vss nfet$245
Xnfet$268_9 m1_n6380_21786# m1_n6380_21786# m1_n6839_21786# m1_n6839_21786# m1_n6282_21430#
+ vss nfet$268
Xnfet$242_78 m1_28010_25858# m1_28634_25662# m1_28371_23922# vss nfet$242
Xnfet$242_67 m1_28492_25858# vss m1_30888_24542# vss nfet$242
Xnfet$242_56 m1_19781_25662# m1_20625_24224# m1_21729_25658# vss nfet$242
Xnfet$242_45 m1_15461_25858# m1_16085_25662# m1_15822_23922# vss nfet$242
Xnfet$242_34 m1_11278_25858# m1_13363_25658# m1_14156_24542# vss nfet$242
Xpfet$228_94 vdd vdd m1_22624_17518# m1_22034_17714# pfet$228
Xpfet$228_83 vdd m1_16538_15778# m1_15921_16080# m1_14641_17836# pfet$228
Xpfet$228_72 vdd m1_20721_15778# m1_20104_16080# m1_18824_17836# pfet$228
Xpfet$228_61 vdd m1_n811_16080# m1_n1278_18030# m1_n2250_17343# pfet$228
Xnfet$242_23 m1_11278_25858# vss m1_11415_25662# vss nfet$242
Xnfet$242_12 m1_7577_25858# vss m1_7522_21786# vss nfet$242
Xpfet$228_50 vdd m1_n1168_15778# m1_n1989_16202# m1_n2250_17343# pfet$228
Xnfet$264_3 m1_n6433_17343# m1_n6172_16202# m1_n6657_17518# vss nfet$264
Xnfet$271_4 m1_n4623_25487# m1_n2567_23922# m1_n3184_24224# vss nfet$271
Xpfet$249_3 vdd m1_n3184_24224# m1_n3651_26174# m1_n4623_25487# pfet$249
Xpfet$227_107 vdd m1_24309_25858# vdd m1_25912_25658# pfet$227
Xnfet$250_9 m1_n7513_20152# vss m1_33790_24346# vss nfet$250
Xnfet$243_8 m1_23486_21590# m1_23486_21590# m1_24973_22513# m1_24973_22513# m1_23945_21586#
+ vss nfet$243
Xpfet$235_9 vdd vdd m1_28624_21786# m1_32675_25947# pfet$235
Xnfet$262_0 m1_4620_20152# m1_4620_20152# m1_2590_19404# m1_2590_19404# m1_3454_20470#
+ vss nfet$262
Xpfet$228_8 vdd vdd m1_9331_15478# sd5 pfet$228
Xpfet$247_0 vdd vdd m1_n7513_20152# m1_35837_22102# pfet$247
Xpfet$254_1 vdd m1_n7186_25858# vdd m1_n6111_25858# pfet$254
Xnfet$241_5 m1_8692_24346# m1_8692_24346# vss vss m1_8174_24542# vss nfet$241
Xnfet$250_12 m1_32675_25947# vss m1_28624_21786# vss nfet$250
Xpfet$233_6 vdd vdd m1_9418_19550# m1_4832_17714# pfet$233
Xpfet$231_3 vdd vdd m1_9418_21590# m1_9288_21786# pfet$231
Xnfet$245_78 m1_14641_17836# m1_15564_15778# m1_14743_16202# vss nfet$245
Xnfet$261_22 m1_15564_15778# m1_15564_15778# m1_15454_18030# m1_15454_18030# m1_15690_17358#
+ vss nfet$261
Xnfet$245_67 m1_17381_17714# vss m1_14482_17343# vss nfet$245
Xnfet$245_56 m1_24287_16080# vss m1_23930_15778# vss nfet$245
Xnfet$245_45 m1_n3064_17714# vss m1_n194_15778# vss nfet$245
Xpfet$227_19 vdd vdd m1_7095_25858# m1_4005_21786# pfet$227
Xnfet$245_34 m1_n2250_17343# vss m1_n2091_17836# vss nfet$245
Xnfet$245_23 m1_5302_17714# vss m1_4832_17714# vss nfet$245
Xnfet$245_12 m1_9485_17714# vss m1_12355_15778# vss nfet$245
Xnfet$261_11 m1_6377_16202# m1_6377_16202# vss vss m1_5859_16398# vss nfet$261
Xnfet$242_79 pd7 vss m1_19839_21786# vss nfet$242
Xnfet$242_68 m1_n7513_20152# vss m1_29607_24346# vss nfet$242
Xnfet$242_57 m1_20126_25858# vss m1_20268_25662# vss nfet$242
Xnfet$242_46 m1_20126_25858# vss m1_18073_21786# vss nfet$242
Xnfet$242_35 m1_15598_25662# m1_15822_23922# m1_16086_24542# vss nfet$242
Xpfet$228_95 vdd vdd m1_21564_17714# m1_22034_17714# pfet$228
Xpfet$228_84 vdd vdd m1_17381_17714# m1_17851_17714# pfet$228
Xpfet$228_73 vdd vdd m1_16538_15778# m1_13668_17714# pfet$228
Xpfet$228_62 vdd vdd m1_23007_17836# m1_22848_17343# pfet$228
Xnfet$242_24 m1_7095_25858# m1_7719_25662# m1_7456_23922# vss nfet$242
Xnfet$242_13 m1_11415_25662# m1_11639_23922# m1_11903_24542# vss nfet$242
Xpfet$228_40 vdd m1_10560_16202# m1_10075_17518# m1_10458_17836# pfet$228
Xpfet$228_51 vdd vdd m1_n1168_15778# m1_n811_16080# pfet$228
Xpfet$230_30 vdd vdd vdd m1_24560_19550# m1_21880_15478# m1_21880_15478# pfet$230
Xnfet$264_4 m1_27031_17343# m1_27292_16202# m1_26807_17518# vss nfet$264
Xnfet$271_5 m1_n4464_25980# m1_n3541_23922# m1_n4362_24346# vss nfet$271
Xpfet$249_4 vdd m1_n2567_23922# m1_n3184_24224# m1_n4464_25980# pfet$249
Xpfet$227_108 vdd vdd m1_25424_24346# m1_n7513_20152# pfet$227
Xnfet$243_9 m1_23356_21786# m1_23356_21786# m1_24973_22513# m1_24973_22513# m1_24577_21586#
+ vss nfet$243
Xnfet$255_0 m1_21456_22513# m1_21456_22513# m1_30256_19792# m1_30256_19792# m1_30492_20470#
+ vss nfet$255
Xnfet$262_1 m1_1103_20152# m1_1103_20152# m1_n927_19404# m1_n927_19404# m1_n63_20470#
+ vss nfet$262
Xpfet$228_9 vdd vdd m1_8172_15778# m1_5302_17714# pfet$228
Xnfet$241_6 m1_8076_24224# m1_8076_24224# m1_7720_24542# m1_7720_24542# m1_8174_24542#
+ vss nfet$241
Xpfet$233_7 vdd vdd m1_11654_20152# m1_5148_15478# pfet$233
Xnfet$250_13 m1_32675_25947# vss m1_32817_25662# vss nfet$250
Xnfet$245_79 m1_15921_16080# vss m1_15564_15778# vss nfet$245
Xnfet$261_23 m1_18926_16202# m1_18926_16202# vss vss m1_18408_16398# vss nfet$261
Xnfet$245_68 m1_18665_17343# m1_18926_16202# m1_18441_17518# vss nfet$245
Xnfet$245_57 m1_22848_17343# m1_24904_15778# m1_24287_16080# vss nfet$245
Xnfet$245_46 m1_22034_17714# vss m1_21564_17714# vss nfet$245
Xnfet$245_24 m1_4832_17714# vss m1_1933_17343# vss nfet$245
Xnfet$245_13 m1_10458_17836# m1_11381_15778# m1_10560_16202# vss nfet$245
Xnfet$245_35 m1_n7513_20152# vss m1_5761_16080# vss nfet$245
Xnfet$261_12 m1_n1168_15778# m1_n1168_15778# m1_n1278_18030# m1_n1278_18030# m1_n1042_17358#
+ vss nfet$261
Xpfet$231_4 vdd vdd m1_8154_21786# m1_7522_21786# pfet$231
Xpfet$228_96 vdd vdd m1_18665_17343# m1_21564_17714# pfet$228
Xpfet$228_85 vdd m1_18926_16202# m1_18441_17518# m1_18824_17836# pfet$228
Xpfet$228_74 vdd vdd m1_14641_17836# m1_14482_17343# pfet$228
Xpfet$228_63 vdd m1_23930_15778# m1_23109_16202# m1_22848_17343# pfet$228
Xpfet$228_30 vdd vdd m1_1933_17343# m1_4832_17714# pfet$228
Xpfet$228_41 vdd vdd m1_10075_17518# m1_9485_17714# pfet$228
Xpfet$228_52 vdd m1_n3064_17714# vdd m1_n1989_16202# pfet$228
Xnfet$242_69 m1_24309_25858# vss m1_26705_24542# vss nfet$242
Xnfet$242_58 m1_20005_23922# vss m1_20625_24224# vss nfet$242
Xnfet$242_47 m1_23964_25662# m1_24188_23922# m1_24452_24542# vss nfet$242
Xnfet$242_36 m1_11760_25858# vss m1_11039_21786# vss nfet$242
Xnfet$242_25 m1_7232_25662# m1_8076_24224# m1_9180_25658# vss nfet$242
Xnfet$242_14 m1_n7513_20152# vss m1_8692_24346# vss nfet$242
Xpfet$230_31 vdd m1_n2543_20130# m1_n2543_20130# m1_20407_19850# m1_19969_19550# m1_19969_19550#
+ pfet$230
Xpfet$230_20 vdd m1_n3822_21786# m1_n3822_21786# m1_14009_19550# m1_9015_17714# m1_9015_17714#
+ pfet$230
Xnfet$264_5 m1_27031_17343# m1_29087_15778# m1_28470_16080# vss nfet$264
Xnfet$271_6 m1_n4464_25980# m1_n3184_24224# m1_n3651_26174# vss nfet$271
Xpfet$249_5 vdd m1_n10572_23922# m1_n10308_24542# m1_n10933_25858# pfet$249
Xpfet$227_109 vdd m1_12259_24224# m1_13363_25658# m1_11278_25858# pfet$227
Xnfet$262_2 m1_n3218_15478# m1_n3218_15478# m1_2590_19404# m1_2590_19404# m1_2822_20470#
+ vss nfet$262
Xnfet$255_1 m1_14422_22513# m1_14422_22513# m1_31535_19792# m1_31535_19792# m1_31771_20470#
+ vss nfet$255
Xnfet$248_0 sd9 vss m1_n7401_15478# vss nfet$248
Xnfet$241_7 m1_9180_25658# m1_9180_25658# vss vss m1_9639_25502# vss nfet$241
Xpfet$233_8 vdd vdd m1_n1133_19550# m1_n7383_17599# pfet$233
Xpfet$252_0 vdd vdd m1_n4485_20152# m1_n3822_20130# pfet$252
Xnfet$261_24 m1_18310_16080# m1_18310_16080# m1_17851_17714# m1_17851_17714# m1_18408_16398#
+ vss nfet$261
Xnfet$245_69 m1_17851_17714# vss m1_17381_17714# vss nfet$245
Xnfet$245_58 m1_23007_17836# m1_23930_15778# m1_23109_16202# vss nfet$245
Xnfet$245_47 m1_22034_17714# vss m1_22624_17518# vss nfet$245
Xnfet$245_25 m1_2092_17836# m1_3372_16080# m1_2905_18030# vss nfet$245
Xnfet$245_14 m1_6116_17343# m1_8172_15778# m1_7555_16080# vss nfet$245
Xnfet$245_36 m1_n3064_17714# vss m1_n2474_17518# vss nfet$245
Xnfet$261_13 m1_n2605_16080# m1_n2605_16080# vss vss m1_n1042_17358# vss nfet$261
Xpfet$231_5 vdd vdd m1_1120_21786# m1_488_21786# pfet$231
Xpfet$228_97 vdd vdd m1_22493_16080# m1_n7513_20152# pfet$228
Xpfet$228_86 vdd m1_19637_18030# vdd m1_18310_16080# pfet$228
Xpfet$228_75 vdd vdd m1_17697_15478# sd3 pfet$228
Xpfet$228_64 vdd vdd m1_23930_15778# m1_24287_16080# pfet$228
Xpfet$228_20 vdd vdd m1_1119_17714# m1_1578_16080# pfet$228
Xpfet$228_31 vdd m1_3372_16080# m1_2905_18030# m1_1933_17343# pfet$228
Xpfet$228_42 vdd m1_11271_18030# vdd m1_9944_16080# pfet$228
Xpfet$228_53 vdd vdd m1_n3218_15478# sd8 pfet$228
Xnfet$242_59 m1_19644_25858# m1_20268_25662# m1_20005_23922# vss nfet$242
Xnfet$242_48 m1_18073_21786# vss m1_23827_25858# vss nfet$242
Xnfet$242_37 m1_11039_21786# vss m1_15461_25858# vss nfet$242
Xnfet$242_26 m1_7095_25858# m1_9180_25658# m1_9973_24542# vss nfet$242
Xnfet$242_15 m1_7232_25662# m1_7456_23922# m1_7720_24542# vss nfet$242
Xpfet$230_32 vdd m1_n2543_20130# m1_n2543_20130# m1_21043_19550# m1_17381_17714# m1_17381_17714#
+ pfet$230
Xpfet$230_21 vdd vdd vdd m1_13373_19850# m1_15171_20152# m1_15171_20152# pfet$230
Xnfet$264_6 m1_27190_17836# m1_28113_15778# m1_27292_16202# vss nfet$264
Xpfet$230_10 vdd vdd vdd m1_9856_19850# m1_11654_20152# m1_11654_20152# pfet$230
Xnfet$271_7 m1_n4623_25487# m1_n4362_24346# m1_n4847_25662# vss nfet$271
Xpfet$249_6 vdd m1_n8848_25658# m1_n8055_24542# m1_n10796_25662# pfet$249
Xnfet$248_1 sd2 vss m1_21880_15478# vss nfet$248
Xnfet$255_2 m1_17939_22513# m1_17939_22513# vss vss m1_31771_20470# vss nfet$255
Xnfet$262_3 m1_8137_20152# m1_8137_20152# m1_6107_19404# m1_6107_19404# m1_6971_20470#
+ vss nfet$262
Xnfet$260_0 fout vss m1_35837_22102# vss nfet$260
Xpfet$233_9 vdd vdd m1_27003_19550# m1_25747_17714# pfet$233
Xnfet$241_8 m1_8692_24346# m1_8692_24346# m1_7577_25858# m1_7577_25858# m1_9639_25502#
+ vss nfet$241
Xpfet$245_0 vdd vdd m1_n7247_17714# m1_n6788_16080# pfet$245
Xpfet$252_1 vdd m1_n4485_21904# vdd m1_9624_19404# pfet$252
Xnfet$245_59 m1_17851_17714# vss m1_20721_15778# vss nfet$245
Xnfet$245_48 m1_18824_17836# m1_20104_16080# m1_19637_18030# vss nfet$245
Xnfet$245_26 m1_5302_17714# vss m1_5892_17518# vss nfet$245
Xnfet$245_15 m1_5302_17714# vss m1_8172_15778# vss nfet$245
Xnfet$245_37 m1_n7513_20152# vss m1_n2605_16080# vss nfet$245
Xpfet$231_6 vdd vdd m1_5901_21590# m1_5771_21786# pfet$231
Xnfet$261_25 m1_14743_16202# m1_14743_16202# vss vss m1_14225_16398# vss nfet$261
Xnfet$261_14 m1_n2605_16080# m1_n2605_16080# m1_n3064_17714# m1_n3064_17714# m1_n2507_16398#
+ vss nfet$261
Xpfet$233_10 vdd vdd m1_29239_20152# m1_26063_15478# pfet$233
Xpfet$228_98 vdd m1_20104_16080# m1_19637_18030# m1_18665_17343# pfet$228
Xpfet$228_87 vdd vdd m1_18310_16080# m1_n7513_20152# pfet$228
Xpfet$228_76 vdd m1_17851_17714# vdd m1_18926_16202# pfet$228
Xpfet$228_65 vdd m1_24904_15778# m1_24287_16080# m1_23007_17836# pfet$228
Xpfet$228_21 vdd vdd m1_965_15478# sd7 pfet$228
Xpfet$228_10 vdd m1_8172_15778# m1_7555_16080# m1_6275_17836# pfet$228
Xpfet$228_32 vdd vdd m1_2905_18030# m1_3015_15778# pfet$228
Xpfet$228_43 vdd vdd m1_11271_18030# m1_11381_15778# pfet$228
Xpfet$228_54 vdd vdd m1_n1278_18030# m1_n1168_15778# pfet$228
Xnfet$242_49 m1_19781_25662# m1_20005_23922# m1_20269_24542# vss nfet$242
Xnfet$242_38 m1_n7513_20152# vss m1_12875_24346# vss nfet$242
Xnfet$242_27 m1_7577_25858# vss m1_7719_25662# vss nfet$242
Xnfet$242_16 m1_4005_21786# vss m1_7095_25858# vss nfet$242
Xnfet$264_7 m1_27190_17836# m1_28470_16080# m1_28003_18030# vss nfet$264
Xpfet$230_33 vdd m1_n3206_20274# m1_n3206_20274# m1_24560_19550# m1_21564_17714# m1_21564_17714#
+ pfet$230
Xpfet$230_22 vdd vdd vdd m1_14009_19550# m1_9331_15478# m1_9331_15478# pfet$230
Xpfet$230_11 vdd vdd vdd m1_10492_19550# m1_5148_15478# m1_5148_15478# pfet$230
Xpfet$249_7 vdd m1_n3541_23922# m1_n4362_24346# m1_n4623_25487# pfet$249
Xnfet$248_2 sd1 vss m1_26063_15478# vss nfet$248
Xnfet$255_3 m1_24973_22513# m1_24973_22513# vss vss m1_30492_20470# vss nfet$255
Xnfet$262_4 m1_965_15478# m1_965_15478# m1_6107_19404# m1_6107_19404# m1_6339_20470#
+ vss nfet$262
Xnfet$241_9 m1_17058_24346# m1_17058_24346# vss vss m1_16540_24542# vss nfet$241
Xnfet$260_1 define m1_35837_22102# vss vss nfet$260
Xpfet$238_0 vdd m1_31535_19792# vdd m1_17939_22513# pfet$238
Xpfet$245_1 vdd m1_n7247_17714# vdd m1_n6172_16202# pfet$245
Xpfet$252_2 vdd m1_n5227_21418# vdd m1_2590_19404# pfet$252
Xnfet$253_0 m1_n290_24224# m1_n290_24224# m1_n646_24542# m1_n646_24542# m1_n192_24542#
+ vss nfet$253
Xpfet$231_7 vdd vdd m1_4637_21786# m1_4005_21786# pfet$231
Xnfet$261_26 m1_14127_16080# m1_14127_16080# m1_13668_17714# m1_13668_17714# m1_14225_16398#
+ vss nfet$261
Xnfet$245_49 m1_21564_17714# vss m1_18665_17343# vss nfet$245
Xnfet$245_27 m1_1119_17714# vss m1_3989_15778# vss nfet$245
Xnfet$245_16 m1_6275_17836# m1_7198_15778# m1_6377_16202# vss nfet$245
Xnfet$245_38 m1_n2250_17343# m1_n1989_16202# m1_n2474_17518# vss nfet$245
Xnfet$261_15 m1_n1989_16202# m1_n1989_16202# vss vss m1_n2507_16398# vss nfet$261
Xpfet$233_11 vdd vdd m1_18688_20152# m1_13514_15478# pfet$233
Xpfet$228_22 vdd vdd m1_3015_15778# m1_3372_16080# pfet$228
Xpfet$228_11 vdd vdd m1_9485_17714# m1_9944_16080# pfet$228
Xpfet$228_33 vdd vdd m1_5892_17518# m1_5302_17714# pfet$228
Xnfet$242_39 pd4 vss m1_9288_21786# vss nfet$242
Xpfet$228_99 vdd m1_23109_16202# m1_22624_17518# m1_23007_17836# pfet$228
Xpfet$228_88 vdd vdd m1_18441_17518# m1_17851_17714# pfet$228
Xpfet$228_77 vdd vdd m1_17851_17714# m1_18310_16080# pfet$228
Xpfet$228_66 vdd vdd m1_24904_15778# m1_22034_17714# pfet$228
Xnfet$242_28 m1_3394_25858# vss m1_4005_21786# vss nfet$242
Xnfet$242_17 m1_11639_23922# vss m1_12259_24224# vss nfet$242
Xpfet$228_44 vdd vdd m1_649_17714# m1_1119_17714# pfet$228
Xpfet$228_55 vdd vdd m1_n2474_17518# m1_n3064_17714# pfet$228
Xpfet$230_34 vdd m1_n3206_20274# m1_n3206_20274# m1_23924_19850# m1_23486_19550# m1_23486_19550#
+ pfet$230
Xpfet$230_23 vdd vdd vdd m1_16890_19850# m1_18688_20152# m1_18688_20152# pfet$230
Xpfet$230_12 vdd m1_6107_19404# m1_6107_19404# m1_6975_19550# m1_649_17714# m1_649_17714#
+ pfet$230
Xnfet$255_4 m1_32818_20470# m1_32818_20470# vss vss m1_34329_20470# vss nfet$255
Xnfet$262_5 m1_5148_15478# m1_5148_15478# m1_9624_19404# m1_9624_19404# m1_9856_20470#
+ vss nfet$262
Xnfet$253_1 m1_814_25658# m1_814_25658# vss vss m1_1273_25502# vss nfet$253
Xpfet$245_2 vdd vdd m1_n5461_18030# m1_n5351_15778# pfet$245
Xnfet$246_0 m1_n1263_21786# vss m1_n1133_21590# vss nfet$246
Xpfet$252_3 vdd vdd m1_n5227_21418# m1_6107_19404# pfet$252
Xpfet$238_1 vdd vdd m1_30256_19792# m1_21456_22513# pfet$238
Xpfet$231_8 vdd vdd m1_2384_21590# m1_2254_21786# pfet$231
Xnfet$261_27 m1_18310_16080# m1_18310_16080# vss vss m1_19873_17358# vss nfet$261
Xnfet$261_16 m1_19747_15778# m1_19747_15778# m1_19637_18030# m1_19637_18030# m1_19873_17358#
+ vss nfet$261
Xnfet$245_28 m1_1933_17343# vss m1_2092_17836# vss nfet$245
Xnfet$245_17 m1_649_17714# vss m1_n2250_17343# vss nfet$245
Xnfet$245_39 m1_n3064_17714# vss m1_n3534_17714# vss nfet$245
Xpfet$250_0 vdd vdd m1_n7320_25516# m1_n7186_25858# pfet$250
Xpfet$233_12 vdd vdd m1_15171_20152# m1_9331_15478# pfet$233
Xnfet$242_29 m1_15943_25858# vss m1_14556_21786# vss nfet$242
Xpfet$228_89 vdd vdd m1_22848_17343# m1_25747_17714# pfet$228
Xpfet$228_78 vdd vdd m1_13514_15478# sd4 pfet$228
Xpfet$228_67 vdd m1_22034_17714# vdd m1_23109_16202# pfet$228
Xnfet$242_18 m1_7095_25858# vss m1_7232_25662# vss nfet$242
Xpfet$228_12 vdd m1_3989_15778# m1_3372_16080# m1_2092_17836# pfet$228
Xpfet$228_23 vdd m1_5302_17714# vdd m1_6377_16202# pfet$228
Xpfet$228_34 vdd vdd m1_5761_16080# m1_n7513_20152# pfet$228
Xpfet$228_45 vdd vdd m1_9944_16080# m1_n7513_20152# pfet$228
Xpfet$228_56 vdd m1_n1278_18030# vdd m1_n2605_16080# pfet$228
Xpfet$230_35 vdd m1_n3822_21786# m1_n3822_21786# m1_13373_19850# m1_12935_19550# m1_12935_19550#
+ pfet$230
Xpfet$230_24 vdd m1_n1927_20274# m1_n1927_20274# m1_16890_19850# m1_16452_19550# m1_16452_19550#
+ pfet$230
Xnfet$276_0 m1_n4485_20152# m1_n6380_21786# vss vss nfet$276
Xpfet$230_13 vdd m1_n927_19404# m1_n927_19404# m1_n695_19850# m1_n1133_19550# m1_n1133_19550#
+ pfet$230
Xnfet$255_5 m1_32818_21586# m1_32818_21586# m1_34093_19792# m1_34093_19792# m1_34329_20470#
+ vss nfet$255
Xnfet$262_6 m1_11654_20152# m1_11654_20152# m1_9624_19404# m1_9624_19404# m1_10488_20470#
+ vss nfet$262
Xnfet$253_2 m1_326_24346# m1_326_24346# m1_n789_25858# m1_n789_25858# m1_1273_25502#
+ vss nfet$253
Xnfet$246_1 m1_11039_21786# vss m1_11671_21786# vss nfet$246
Xpfet$238_2 vdd m1_30256_19792# vdd m1_24973_22513# pfet$238
Xpfet$245_3 vdd m1_n5461_18030# vdd m1_n6788_16080# pfet$245
Xpfet$252_4 vdd vdd m1_n4485_21904# m1_n3822_21786# pfet$252
Xpfet$243_0 vdd vdd fout m1_34093_22102# pfet$243
Xpfet$231_9 vdd vdd m1_22222_21786# m1_21590_21786# pfet$231
Xnfet$261_17 m1_22493_16080# m1_22493_16080# vss vss m1_24056_17358# vss nfet$261
Xnfet$245_29 m1_3372_16080# vss m1_3015_15778# vss nfet$245
Xnfet$245_18 m1_1119_17714# vss m1_649_17714# vss nfet$245
Xpfet$250_1 vdd vdd m1_n6111_25858# m1_n6856_24542# pfet$250
Xpfet$233_13 vdd vdd m1_16452_19550# m1_13198_17714# pfet$233
Xpfet$228_79 vdd m1_15564_15778# m1_14743_16202# m1_14482_17343# pfet$228
Xpfet$228_68 vdd vdd m1_22034_17714# m1_22493_16080# pfet$228
Xpfet$228_13 vdd vdd m1_5148_15478# sd6 pfet$228
Xpfet$228_24 vdd m1_6377_16202# m1_5892_17518# m1_6275_17836# pfet$228
Xpfet$228_35 vdd vdd m1_9015_17714# m1_9485_17714# pfet$228
Xpfet$228_46 vdd vdd m1_n2250_17343# m1_649_17714# pfet$228
Xpfet$228_57 vdd m1_n1989_16202# m1_n2474_17518# m1_n2091_17836# pfet$228
Xnfet$242_19 m1_7456_23922# vss m1_8076_24224# vss nfet$242
Xpfet$230_25 vdd vdd vdd m1_17526_19550# m1_13514_15478# m1_13514_15478# pfet$230
Xpfet$230_14 vdd m1_n927_19404# m1_n927_19404# m1_n59_19550# m1_n7383_17599# m1_n7383_17599#
+ pfet$230
Xnfet$276_1 m1_n5227_20152# vss m1_n6380_21786# vss nfet$276
Xnfet$269_0 m1_n8625_26174# vss m1_n8055_24542# vss nfet$269
Xnfet$262_7 m1_n7401_15478# m1_n7401_15478# m1_n927_19404# m1_n927_19404# m1_n695_20470#
+ vss nfet$262
Xnfet$255_6 m1_354_22513# m1_354_22513# m1_31535_22102# m1_31535_22102# m1_31771_21430#
+ vss nfet$255
Xnfet$253_3 m1_326_24346# m1_326_24346# vss vss m1_n192_24542# vss nfet$253
Xnfet$246_2 m1_12805_21786# vss m1_12935_21590# vss nfet$246
Xpfet$238_3 vdd vdd m1_34843_21786# m1_34093_19792# pfet$238
Xpfet$245_4 vdd vdd m1_26217_17714# m1_26676_16080# pfet$245
Xpfet$252_5 vdd m1_n6839_21786# vdd m1_n5764_21786# pfet$252
Xnfet$261_18 m1_23930_15778# m1_23930_15778# m1_23820_18030# m1_23820_18030# m1_24056_17358#
+ vss nfet$261
Xnfet$245_19 m1_n7513_20152# vss m1_1578_16080# vss nfet$245
Xnfet$251_0 m1_n1134_25662# m1_n910_23922# m1_n646_24542# vss nfet$251
Xpfet$236_0 vdd vdd m1_n646_24542# m1_n290_24224# pfet$236
Xpfet$233_14 vdd vdd m1_23486_19550# m1_21564_17714# pfet$233
Xpfet$228_69 vdd vdd m1_20721_15778# m1_17851_17714# pfet$228
Xpfet$228_14 vdd vdd m1_2092_17836# m1_1933_17343# pfet$228
Xpfet$228_25 vdd vdd m1_1709_17518# m1_1119_17714# pfet$228
Xpfet$228_36 vdd vdd m1_6116_17343# m1_9015_17714# pfet$228
Xpfet$228_47 vdd m1_11738_16080# m1_11271_18030# m1_10299_17343# pfet$228
Xpfet$228_58 vdd vdd m1_n3534_17714# m1_n3064_17714# pfet$228
Xpfet$230_26 vdd m1_n1927_20274# m1_n1927_20274# m1_17526_19550# m1_13198_17714# m1_13198_17714#
+ pfet$230
Xpfet$230_15 vdd vdd vdd m1_n59_19550# m1_n7401_15478# m1_n7401_15478# pfet$230
Xnfet$269_1 m1_n8625_26174# vss m1_n7082_23622# vss nfet$269
Xnfet$255_7 m1_3871_22513# m1_3871_22513# vss vss m1_31771_21430# vss nfet$255
Xnfet$262_8 m1_26063_15478# m1_26063_15478# m1_n3822_20130# m1_n3822_20130# m1_27441_20470#
+ vss nfet$262
Xnfet$253_4 m1_33174_24224# m1_33174_24224# m1_32818_24542# m1_32818_24542# m1_33272_24542#
+ vss nfet$253
Xnfet$246_3 m1_9288_21786# vss m1_9418_21590# vss nfet$246
Xpfet$238_4 vdd m1_34093_19792# vdd m1_32818_20470# pfet$238
Xpfet$245_5 vdd m1_26217_17714# vdd m1_27292_16202# pfet$245
Xpfet$252_6 vdd vdd m1_n6973_21481# m1_n6839_21786# pfet$252
Xnfet$244_0 m1_n3534_17714# m1_n3534_17714# vss vss m1_3454_20470# vss nfet$244
Xnfet$251_1 m1_n1271_25858# m1_n647_25662# m1_n910_23922# vss nfet$251
Xnfet$261_19 m1_23109_16202# m1_23109_16202# vss vss m1_22591_16398# vss nfet$261
Xpfet$236_1 vdd m1_n789_25858# vdd m1_814_25658# pfet$236
Xpfet$229_0 vdd vdd vdd m1_n674_22102# m1_n1133_21590# m1_n1133_21590# pfet$229
Xpfet$233_15 vdd vdd m1_22205_20152# m1_17697_15478# pfet$233
Xpfet$228_15 vdd vdd m1_5302_17714# m1_5761_16080# pfet$228
Xpfet$228_26 vdd vdd m1_4832_17714# m1_5302_17714# pfet$228
Xpfet$228_37 vdd m1_7555_16080# m1_7088_18030# m1_6116_17343# pfet$228
Xpfet$228_48 vdd vdd m1_n3064_17714# m1_n2605_16080# pfet$228
Xpfet$228_59 vdd vdd m1_n2605_16080# m1_n7513_20152# pfet$228
Xpfet$230_27 vdd vdd vdd m1_20407_19850# m1_22205_20152# m1_22205_20152# pfet$230
Xpfet$230_16 vdd vdd vdd m1_28077_19550# m1_26063_15478# m1_26063_15478# pfet$230
Xnfet$269_2 vss vss m1_n9336_24346# vss nfet$269
Xnfet$262_9 m1_29239_20152# m1_29239_20152# m1_n3822_20130# m1_n3822_20130# m1_28073_20470#
+ vss nfet$262
Xpfet$259_0 vdd vdd m1_n8145_21908# m1_n6839_20152# pfet$259
Xnfet$274_0 m1_n4485_21904# m1_n5764_21786# vss vss nfet$274
Xnfet$253_5 m1_33790_24346# m1_33790_24346# vss vss m1_33272_24542# vss nfet$253
Xpfet$245_6 vdd vdd m1_28003_18030# m1_28113_15778# pfet$245
Xpfet$238_5 vdd vdd m1_34093_19792# m1_32818_21586# pfet$238
Xpfet$252_7 vdd vdd m1_n6839_21786# m1_n6380_21786# pfet$252
Xnfet$246_4 m1_7522_21786# vss m1_8154_21786# vss nfet$246
Xnfet$244_1 m1_2384_19550# m1_2384_19550# vss vss m1_2822_20470# vss nfet$244
Xnfet$251_2 m1_n1271_25858# m1_814_25658# m1_1607_24542# vss nfet$251
Xpfet$236_2 vdd vdd m1_n789_25858# m1_326_24346# pfet$236
Xpfet$229_1 vdd m1_7388_22513# m1_7388_22513# m1_6988_22402# m1_7522_21786# m1_7522_21786#
+ pfet$229
Xpfet$233_16 vdd vdd m1_19969_19550# m1_17381_17714# pfet$233
Xpfet$241_0 vdd m1_34093_22102# vdd m1_28490_22513# pfet$241
Xpfet$228_16 vdd vdd m1_3989_15778# m1_1119_17714# pfet$228
Xpfet$228_27 vdd m1_2194_16202# m1_1709_17518# m1_2092_17836# pfet$228
Xpfet$228_38 vdd vdd m1_7088_18030# m1_7198_15778# pfet$228
Xpfet$228_49 vdd m1_n194_15778# m1_n811_16080# m1_n2091_17836# pfet$228
Xpfet$230_28 vdd vdd vdd m1_21043_19550# m1_17697_15478# m1_17697_15478# pfet$230
Xpfet$230_17 vdd m1_n3822_20130# m1_n3822_20130# m1_28077_19550# m1_25747_17714# m1_25747_17714#
+ pfet$230
Xnfet$269_3 fin vss m1_n10933_25858# vss nfet$269
Xnfet$243_10 m1_19839_21786# m1_19839_21786# m1_21456_22513# m1_21456_22513# m1_21060_21586#
+ vss nfet$243
Xnfet$274_1 m1_n5227_21418# vss m1_n5764_21786# vss nfet$274
Xnfet$267_0 m1_n7082_23622# m1_n6856_24542# vss vss nfet$267
Xnfet$253_6 m1_33790_24346# m1_33790_24346# m1_32675_25947# m1_32675_25947# m1_34737_25502#
+ vss nfet$253
Xpfet$245_7 vdd m1_28003_18030# vdd m1_26676_16080# pfet$245
Xnfet$246_5 m1_488_21786# vss m1_1120_21786# vss nfet$246
Xpfet$238_6 vdd vdd m1_31535_19792# m1_14422_22513# pfet$238
Xnfet$251_3 m1_n1134_25662# m1_n290_24224# m1_814_25658# vss nfet$251
Xpfet$236_3 vdd m1_n646_24542# vdd m1_326_24346# pfet$236
Xnfet$244_2 m1_5901_19550# m1_5901_19550# vss vss m1_6339_20470# vss nfet$244
Xpfet$229_2 vdd m1_7388_22513# m1_7388_22513# m1_6360_22102# m1_8154_21786# m1_8154_21786#
+ pfet$229
Xpfet$233_17 vdd vdd m1_25722_20152# m1_21880_15478# pfet$233
Xpfet$241_1 vdd vdd m1_34093_22102# m1_34843_21786# pfet$241
Xnfet$246_10 m1_21590_21786# vss m1_22222_21786# vss nfet$246
Xpfet$234_0 vdd vdd m1_n7401_15478# sd9 pfet$234
Xpfet$228_17 vdd vdd m1_n2091_17836# m1_n2250_17343# pfet$228
Xpfet$228_28 vdd m1_2905_18030# vdd m1_1578_16080# pfet$228
Xpfet$228_39 vdd m1_7088_18030# vdd m1_5761_16080# pfet$228
Xpfet$230_29 vdd vdd vdd m1_23924_19850# m1_25722_20152# m1_25722_20152# pfet$230
Xpfet$230_18 vdd vdd vdd m1_27441_19850# m1_29239_20152# m1_29239_20152# pfet$230
Xnfet$269_4 m1_n10572_23922# vss m1_n9952_24224# vss nfet$269
Xnfet$243_11 m1_19969_21590# m1_19969_21590# m1_21456_22513# m1_21456_22513# m1_20428_21586#
+ vss nfet$243
Xnfet$274_2 m1_n6839_21786# vss m1_n6973_21481# vss nfet$274
Xnfet$267_1 m1_n8283_19850# vss m1_n6856_24542# vss nfet$267
Xnfet$254_10 m1_21590_21786# m1_21590_21786# vss vss m1_20428_21586# vss nfet$254
Xnfet$253_7 m1_34278_25658# m1_34278_25658# vss vss m1_34737_25502# vss nfet$253
Xnfet$246_6 m1_5771_21786# vss m1_5901_21590# vss nfet$246
Xpfet$238_7 vdd vdd m1_31535_22102# m1_354_22513# pfet$238
Xnfet$249_10 m1_26217_17714# vss m1_29087_15778# vss nfet$249
Xpfet$236_4 vdd vdd m1_32675_25947# m1_33790_24346# pfet$236
Xnfet$251_4 m1_32193_25858# m1_34278_25658# m1_35071_24542# vss nfet$251
Xnfet$244_3 m1_4832_17714# m1_4832_17714# vss vss m1_10488_20470# vss nfet$244
Xpfet$229_3 vdd m1_9645_21447# m1_9645_21447# m1_10505_22402# m1_11039_21786# m1_11039_21786#
+ pfet$229
Xnfet$242_0 m1_3394_25858# vss m1_5790_24542# vss nfet$242
Xpfet$241_2 vdd vdd m1_30256_22102# m1_7388_22513# pfet$241
Xnfet$246_11 m1_18073_21786# vss m1_18705_21786# vss nfet$246
Xpfet$234_1 vdd vdd m1_21880_15478# sd2 pfet$234
Xpfet$227_0 vdd vdd m1_3049_25662# m1_2912_25858# pfet$227
Xnfet$262_10 m1_9331_15478# m1_9331_15478# m1_n3822_21786# m1_n3822_21786# m1_13373_20470#
+ vss nfet$262
Xpfet$228_18 vdd m1_1119_17714# vdd m1_2194_16202# pfet$228
Xpfet$228_29 vdd vdd m1_1578_16080# m1_n7513_20152# pfet$228
Xpfet$230_19 vdd m1_n3822_20130# m1_n3822_20130# m1_27441_19850# m1_27003_19550# m1_27003_19550#
+ pfet$230
Xnfet$269_5 m1_n10933_25858# vss m1_n10796_25662# vss nfet$269
Xnfet$243_12 m1_16322_21786# m1_16322_21786# m1_17939_22513# m1_17939_22513# m1_17543_21586#
+ vss nfet$243
Xnfet$254_11 m1_22222_21786# m1_22222_21786# vss vss m1_21060_21586# vss nfet$254
Xnfet$246_7 m1_4005_21786# vss m1_4637_21786# vss nfet$246
Xnfet$272_0 m1_n7186_25858# vss m1_n7320_25516# vss nfet$272
Xnfet$249_11 m1_27031_17343# vss m1_27190_17836# vss nfet$249
Xpfet$257_0 vdd vdd m1_n5227_20152# m1_n2543_20130# pfet$257
Xnfet$251_5 m1_32330_25662# m1_33174_24224# m1_34278_25658# vss nfet$251
Xnfet$244_4 m1_9418_19550# m1_9418_19550# vss vss m1_9856_20470# vss nfet$244
Xpfet$236_5 vdd m1_32675_25947# vdd m1_34278_25658# pfet$236
Xpfet$229_4 vdd vdd vdd m1_9877_22102# m1_9418_21590# m1_9418_21590# pfet$229
Xpfet$234_2 vdd vdd m1_26063_15478# sd1 pfet$234
Xpfet$241_3 vdd m1_31535_22102# vdd m1_3871_22513# pfet$241
Xpfet$227_1 vdd m1_3536_25662# m1_3273_23922# m1_3049_25662# pfet$227
Xnfet$242_1 m1_2912_25858# m1_4997_25658# m1_5790_24542# vss nfet$242
Xnfet$246_12 m1_14556_21786# vss m1_15188_21786# vss nfet$246
Xnfet$262_11 m1_15171_20152# m1_15171_20152# m1_n3822_21786# m1_n3822_21786# m1_14005_20470#
+ vss nfet$262
Xpfet$228_19 vdd m1_3015_15778# m1_2194_16202# m1_1933_17343# pfet$228
Xnfet$269_6 m1_n10452_25858# vss m1_n10309_25662# vss nfet$269
Xnfet$243_13 m1_16452_21590# m1_16452_21590# m1_17939_22513# m1_17939_22513# m1_16911_21586#
+ vss nfet$243
Xnfet$254_12 m1_18073_21786# m1_18073_21786# vss vss m1_16911_21586# vss nfet$254
Xnfet$246_8 m1_2254_21786# vss m1_2384_21590# vss nfet$246
Xnfet$265_0 m1_n5351_15778# m1_n5351_15778# m1_n5461_18030# m1_n5461_18030# m1_n5225_17358#
+ vss nfet$265
Xnfet$272_1 m1_n6856_24542# vss m1_n6111_25858# vss nfet$272
Xnfet$249_12 m1_28470_16080# vss m1_28113_15778# vss nfet$249
Xpfet$257_1 vdd m1_n4485_20152# vdd m1_n3206_20274# pfet$257
Xnfet$251_6 m1_32193_25858# m1_32817_25662# m1_32554_23922# vss nfet$251
Xnfet$244_5 m1_649_17714# m1_649_17714# vss vss m1_6971_20470# vss nfet$244
Xpfet$236_6 vdd vdd m1_32818_24542# m1_33174_24224# pfet$236
Xpfet$229_5 vdd m1_9645_21447# m1_9645_21447# m1_9877_22102# m1_11671_21786# m1_11671_21786#
+ pfet$229
Xpfet$241_4 vdd m1_30256_22102# vdd m1_9645_21447# pfet$241
Xnfet$242_2 m1_n7513_20152# vss m1_4509_24346# vss nfet$242
Xnfet$246_13 m1_16322_21786# vss m1_16452_21590# vss nfet$246
Xnfet$262_12 m1_18688_20152# m1_18688_20152# m1_n1927_20274# m1_n1927_20274# m1_17522_20470#
+ vss nfet$262
Xpfet$227_2 vdd vdd m1_3394_25858# m1_4509_24346# pfet$227
Xpfet$232_0 vdd vdd m1_n6274_17836# m1_n6433_17343# pfet$232
Xnfet$269_7 m1_n7320_25516# vss m1_n2567_23922# vss nfet$269
Xpfet$229_30 vdd vdd vdd m1_17539_22402# m1_16322_21786# m1_16322_21786# pfet$229
Xnfet$243_14 m1_12805_21786# m1_12805_21786# m1_14422_22513# m1_14422_22513# m1_14026_21586#
+ vss nfet$243
Xnfet$254_13 m1_18705_21786# m1_18705_21786# vss vss m1_17543_21586# vss nfet$254
Xnfet$246_9 m1_23356_21786# vss m1_23486_21590# vss nfet$246
Xnfet$258_0 m1_34093_19792# vss m1_34843_21786# vss nfet$258
Xnfet$265_1 m1_n6788_16080# m1_n6788_16080# vss vss m1_n5225_17358# vss nfet$265
Xnfet$249_13 m1_26217_17714# vss m1_25747_17714# vss nfet$249
Xpfet$257_2 vdd m1_n5227_20152# vdd m1_n1927_20274# pfet$257
Xnfet$251_7 m1_32330_25662# m1_32554_23922# m1_32818_24542# vss nfet$251
Xnfet$244_6 m1_n1133_19550# m1_n1133_19550# vss vss m1_n695_20470# vss nfet$244
Xpfet$236_7 vdd m1_32818_24542# vdd m1_33790_24346# pfet$236
Xpfet$229_6 vdd vdd vdd m1_10505_22402# m1_9288_21786# m1_9288_21786# pfet$229
Xnfet$242_3 m1_488_21786# vss m1_2912_25858# vss nfet$242
Xnfet$246_14 m1_19839_21786# vss m1_19969_21590# vss nfet$246
Xnfet$262_13 m1_13514_15478# m1_13514_15478# m1_n1927_20274# m1_n1927_20274# m1_16890_20470#
+ vss nfet$262
Xpfet$227_3 vdd m1_3394_25858# vdd m1_4997_25658# pfet$227
Xpfet$232_1 vdd vdd m1_n4377_15778# m1_n7247_17714# pfet$232
Xnfet$269_8 m1_n4623_25487# vss m1_n4464_25980# vss nfet$269
Xpfet$229_31 vdd vdd vdd m1_27462_22102# m1_27003_21590# m1_27003_21590# pfet$229
Xpfet$229_20 vdd vdd vdd m1_20428_22102# m1_19969_21590# m1_19969_21590# pfet$229
Xnfet$243_15 m1_26873_21786# m1_26873_21786# m1_28490_22513# m1_28490_22513# m1_28094_21586#
+ vss nfet$243
Xpfet$231_10 vdd vdd m1_23486_21590# m1_23356_21786# pfet$231
Xnfet$254_14 m1_15188_21786# m1_15188_21786# vss vss m1_14026_21586# vss nfet$254
Xnfet$258_1 m1_30256_19792# vss m1_32818_20470# vss nfet$258
Xnfet$265_2 m1_n6788_16080# m1_n6788_16080# m1_n7247_17714# m1_n7247_17714# m1_n6690_16398#
+ vss nfet$265
Xpfet$257_3 vdd m1_n6839_20152# vdd m1_n927_19404# pfet$257
Xnfet$244_7 m1_n7383_17599# m1_n7383_17599# vss vss m1_n63_20470# vss nfet$244
Xnfet$270_0 m1_n9952_24224# m1_n9952_24224# m1_n10308_24542# m1_n10308_24542# m1_n9854_24542#
+ vss nfet$270
Xpfet$229_7 vdd m1_354_22513# m1_354_22513# m1_n674_22102# m1_1120_21786# m1_1120_21786#
+ pfet$229
Xpfet$255_0 vdd vdd vdd m1_n8047_19550# m1_n7513_20152# m1_n7513_20152# pfet$255
Xnfet$242_4 m1_2912_25858# vss m1_3049_25662# vss nfet$242
Xnfet$246_15 m1_28624_21786# vss m1_29256_21786# vss nfet$246
Xnfet$262_14 m1_22205_20152# m1_22205_20152# m1_n2543_20130# m1_n2543_20130# m1_21039_20470#
+ vss nfet$262
Xpfet$227_4 vdd vdd m1_3893_24224# m1_3273_23922# pfet$227
Xpfet$232_2 vdd vdd m1_n5351_15778# m1_n4994_16080# pfet$232
Xnfet$269_9 m1_n3184_24224# vss m1_n3541_23922# vss nfet$269
Xpfet$229_32 vdd m1_28490_22513# m1_28490_22513# m1_28090_22402# m1_28624_21786# m1_28624_21786#
+ pfet$229
Xpfet$229_21 vdd vdd vdd m1_21056_22402# m1_19839_21786# m1_19839_21786# pfet$229
Xpfet$229_10 vdd m1_3871_22513# m1_3871_22513# m1_2843_22102# m1_4637_21786# m1_4637_21786#
+ pfet$229
Xnfet$243_16 m1_27003_21590# m1_27003_21590# m1_28490_22513# m1_28490_22513# m1_27462_21586#
+ vss nfet$243
Xpfet$231_11 vdd vdd m1_18705_21786# m1_18073_21786# pfet$231
Xnfet$254_15 m1_14556_21786# m1_14556_21786# vss vss m1_13394_21586# vss nfet$254
Xnfet$258_2 m1_31535_19792# m1_32818_20470# vss vss nfet$258
Xnfet$265_3 m1_n6172_16202# m1_n6172_16202# vss vss m1_n6690_16398# vss nfet$265
Xpfet$257_4 vdd vdd m1_n6839_20152# m1_n6973_21481# pfet$257
Xnfet$263_0 m1_35837_22102# vss m1_n7513_20152# vss nfet$263
Xnfet$244_8 m1_27003_19550# m1_27003_19550# vss vss m1_27441_20470# vss nfet$244
Xnfet$270_1 m1_n9336_24346# m1_n9336_24346# m1_n8625_26174# m1_n8625_26174# m1_n8389_25502#
+ vss nfet$270
Xpfet$229_8 vdd vdd vdd m1_6360_22102# m1_5901_21590# m1_5901_21590# pfet$229
Xpfet$255_1 vdd m1_n8283_19850# m1_n8283_19850# m1_n8047_19550# m1_n8283_20611# m1_n8283_20611#
+ pfet$255
Xpfet$248_0 vdd vdd vdd m1_n6624_23622# m1_n7082_23622# m1_n7082_23622# pfet$248
Xnfet$242_5 m1_2912_25858# m1_3536_25662# m1_3273_23922# vss nfet$242
Xnfet$246_16 m1_26873_21786# vss m1_27003_21590# vss nfet$246
Xpfet$227_5 vdd m1_3893_24224# m1_4997_25658# m1_2912_25858# pfet$227
Xnfet$262_15 m1_17697_15478# m1_17697_15478# m1_n2543_20130# m1_n2543_20130# m1_20407_20470#
+ vss nfet$262
Xpfet$232_3 vdd vdd m1_n6657_17518# m1_n7247_17714# pfet$232
Xpfet$228_110 vdd vdd m1_10458_17836# m1_10299_17343# pfet$228
Xpfet$229_33 vdd m1_28490_22513# m1_28490_22513# m1_27462_22102# m1_29256_21786# m1_29256_21786#
+ pfet$229
Xpfet$229_22 vdd m1_21456_22513# m1_21456_22513# m1_20428_22102# m1_22222_21786# m1_22222_21786#
+ pfet$229
Xpfet$229_11 vdd vdd vdd m1_2843_22102# m1_2384_21590# m1_2384_21590# pfet$229
Xnfet$243_17 m1_12935_21590# m1_12935_21590# m1_14422_22513# m1_14422_22513# m1_13394_21586#
+ vss nfet$243
Xpfet$230_0 vdd m1_2590_19404# m1_2590_19404# m1_3458_19550# m1_n3534_17714# m1_n3534_17714#
+ pfet$230
Xpfet$231_12 vdd vdd m1_16452_21590# m1_16322_21786# pfet$231
Xnfet$254_16 m1_28624_21786# m1_28624_21786# vss vss m1_27462_21586# vss nfet$254
Xnfet$258_3 m1_30256_22102# vss m1_32818_21586# vss nfet$258
Xnfet$265_4 m1_28113_15778# m1_28113_15778# m1_28003_18030# m1_28003_18030# m1_28239_17358#
+ vss nfet$265
Xnfet$244_9 m1_25747_17714# m1_25747_17714# vss vss m1_28073_20470# vss nfet$244
Xnfet$256_0 m1_34843_21786# m1_34843_21786# m1_34093_22102# m1_34093_22102# m1_34329_21430#
+ vss nfet$256
Xpfet$255_2 vdd m1_n8283_20611# m1_n8283_20611# m1_n8047_22344# m1_n8145_21908# m1_n8145_21908#
+ pfet$255
Xnfet$270_2 m1_n8848_25658# m1_n8848_25658# vss vss m1_n8389_25502# vss nfet$270
Xpfet$253_10 vdd vdd m1_n10933_25858# fin pfet$253
Xpfet$248_1 vdd m1_n6856_24542# m1_n6856_24542# m1_n6624_23622# m1_n8283_19850# m1_n8283_19850#
+ pfet$248
Xpfet$229_9 vdd m1_3871_22513# m1_3871_22513# m1_3471_22402# m1_4005_21786# m1_4005_21786#
+ pfet$229
Xpfet$227_6 vdd vdd m1_3536_25662# m1_3394_25858# pfet$227
Xnfet$242_6 m1_3049_25662# m1_3893_24224# m1_4997_25658# vss nfet$242
Xnfet$246_17 m1_25107_21786# vss m1_25739_21786# vss nfet$246
Xnfet$262_16 m1_25722_20152# m1_25722_20152# m1_n3206_20274# m1_n3206_20274# m1_24556_20470#
+ vss nfet$262
Xpfet$232_4 vdd vdd m1_n6433_17343# m1_n3534_17714# pfet$232
Xpfet$229_12 vdd vdd vdd m1_3471_22402# m1_2254_21786# m1_2254_21786# pfet$229
Xpfet$229_34 vdd vdd vdd m1_28090_22402# m1_26873_21786# m1_26873_21786# pfet$229
Xpfet$229_23 vdd vdd vdd m1_23945_22102# m1_23486_21590# m1_23486_21590# pfet$229
Xpfet$228_100 vdd vdd m1_23820_18030# m1_23930_15778# pfet$228
Xpfet$230_1 vdd vdd vdd m1_2822_19850# m1_4620_20152# m1_4620_20152# pfet$230
Xpfet$231_13 vdd vdd m1_15188_21786# m1_14556_21786# pfet$231
Xnfet$254_17 m1_29256_21786# m1_29256_21786# vss vss m1_28094_21586# vss nfet$254
Xnfet$265_5 m1_26676_16080# m1_26676_16080# vss vss m1_28239_17358# vss nfet$265
Xnfet$256_1 m1_28490_22513# m1_28490_22513# vss vss m1_34329_21430# vss nfet$256
Xnfet$249_0 m1_n3534_17714# vss m1_n6433_17343# vss nfet$249
Xnfet$270_3 m1_n9336_24346# m1_n9336_24346# vss vss m1_n9854_24542# vss nfet$270
Xpfet$253_11 vdd vdd m1_n9336_24346# vss pfet$253
Xpfet$255_3 vdd vdd vdd m1_n8047_22344# m1_n8283_19850# m1_n8283_19850# pfet$255
Xnfet$242_7 m1_3049_25662# m1_3273_23922# m1_3537_24542# vss nfet$242
Xnfet$262_17 m1_21880_15478# m1_21880_15478# m1_n3206_20274# m1_n3206_20274# m1_23924_20470#
+ vss nfet$262
Xpfet$227_7 vdd vdd m1_7232_25662# m1_7095_25858# pfet$227
Xpfet$253_0 vdd vdd m1_n10796_25662# m1_n10933_25858# pfet$253
Xpfet$232_5 vdd vdd m1_n6788_16080# m1_n7513_20152# pfet$232
Xpfet$229_35 vdd vdd vdd m1_13394_22102# m1_12935_21590# m1_12935_21590# pfet$229
Xpfet$229_24 vdd m1_17939_22513# m1_17939_22513# m1_16911_22102# m1_18705_21786# m1_18705_21786#
+ pfet$229
Xpfet$228_101 vdd vdd m1_19637_18030# m1_19747_15778# pfet$228
Xpfet$229_13 vdd vdd vdd m1_6988_22402# m1_5771_21786# m1_5771_21786# pfet$229
Xpfet$230_2 vdd m1_2590_19404# m1_2590_19404# m1_2822_19850# m1_2384_19550# m1_2384_19550#
+ pfet$230
Xpfet$231_14 vdd vdd m1_19969_21590# m1_19839_21786# pfet$231
Xnfet$265_6 m1_27292_16202# m1_27292_16202# vss vss m1_26774_16398# vss nfet$265
Xnfet$256_2 m1_9645_21447# m1_9645_21447# vss vss m1_30492_21430# vss nfet$256
Xnfet$249_1 m1_n7513_20152# vss m1_n6788_16080# vss nfet$249
Xnfet$270_4 m1_n4978_24224# m1_n4978_24224# m1_n10452_25858# m1_n10452_25858# m1_n4880_24542#
+ vss nfet$270
Xpfet$253_12 vdd vdd m1_n7082_23622# m1_n8625_26174# pfet$253
Xpfet$227_90 vdd vdd m1_24309_25858# m1_25424_24346# pfet$227
Xnfet$242_8 m1_3394_25858# vss m1_3536_25662# vss nfet$242
Xpfet$227_8 vdd vdd m1_8076_24224# m1_7456_23922# pfet$227
Xnfet$261_0 m1_7198_15778# m1_7198_15778# m1_7088_18030# m1_7088_18030# m1_7324_17358#
+ vss nfet$261
Xpfet$246_0 vdd m1_n4377_15778# m1_n4994_16080# m1_n6274_17836# pfet$246
Xpfet$253_1 vdd vdd m1_n10309_25662# m1_n10452_25858# pfet$253
Xpfet$232_6 vdd vdd m1_n7383_17599# m1_n7247_17714# pfet$232
Xpfet$229_25 vdd m1_17939_22513# m1_17939_22513# m1_17539_22402# m1_18073_21786# m1_18073_21786#
+ pfet$229
Xpfet$228_102 vdd vdd m1_13198_17714# m1_13668_17714# pfet$228
Xpfet$229_14 vdd vdd vdd m1_n46_22402# m1_n1263_21786# m1_n1263_21786# pfet$229
Xpfet$230_3 vdd vdd vdd m1_3458_19550# m1_n3218_15478# m1_n3218_15478# pfet$230
Xpfet$231_15 vdd vdd m1_27003_21590# m1_26873_21786# pfet$231
Xnfet$265_7 m1_26676_16080# m1_26676_16080# m1_26217_17714# m1_26217_17714# m1_26774_16398#
+ vss nfet$265
Xnfet$256_3 m1_7388_22513# m1_7388_22513# m1_30256_22102# m1_30256_22102# m1_30492_21430#
+ vss nfet$256
Xnfet$249_2 m1_n4994_16080# vss m1_n5351_15778# vss nfet$249
Xnfet$270_5 m1_n4362_24346# m1_n4362_24346# vss vss m1_n4880_24542# vss nfet$270
Xpfet$253_13 vdd vdd m1_n8055_24542# m1_n8625_26174# pfet$253
Xpfet$227_91 vdd vdd m1_23356_21786# pd8 pfet$227
Xpfet$227_80 vdd vdd m1_17058_24346# m1_n7513_20152# pfet$227
Xnfet$241_20 m1_21241_24346# m1_21241_24346# m1_20126_25858# m1_20126_25858# m1_22188_25502#
+ vss nfet$241
Xnfet$242_9 m1_3273_23922# vss m1_3893_24224# vss nfet$242
Xpfet$227_9 vdd m1_7719_25662# m1_7456_23922# m1_7232_25662# pfet$227
Xnfet$261_1 m1_5761_16080# m1_5761_16080# vss vss m1_7324_17358# vss nfet$261
Xnfet$254_0 m1_11039_21786# m1_11039_21786# vss vss m1_9877_21586# vss nfet$254
Xpfet$246_1 vdd m1_n5351_15778# m1_n6172_16202# m1_n6433_17343# pfet$246
Xpfet$253_2 vdd vdd m1_n9952_24224# m1_n10572_23922# pfet$253
Xpfet$239_0 vdd m1_n647_25662# m1_n910_23922# m1_n1134_25662# pfet$239
Xpfet$232_7 vdd vdd m1_27190_17836# m1_27031_17343# pfet$232
Xpfet$229_26 vdd vdd vdd m1_16911_22102# m1_16452_21590# m1_16452_21590# pfet$229
Xpfet$228_103 vdd m1_14743_16202# m1_14258_17518# m1_14641_17836# pfet$228
Xpfet$229_15 vdd m1_354_22513# m1_354_22513# m1_n46_22402# m1_488_21786# m1_488_21786#
+ pfet$229
Xpfet$230_4 vdd m1_6107_19404# m1_6107_19404# m1_6339_19850# m1_5901_19550# m1_5901_19550#
+ pfet$230
Xpfet$231_16 vdd vdd m1_29256_21786# m1_28624_21786# pfet$231
Xnfet$270_6 m1_n4978_24224# m1_n4978_24224# vss vss m1_n3415_25502# vss nfet$270
Xpfet$227_92 vdd vdd m1_28492_25858# m1_29607_24346# pfet$227
Xpfet$227_81 vdd vdd m1_18339_24542# m1_15943_25858# pfet$227
Xpfet$227_70 vdd vdd m1_14156_24542# m1_11760_25858# pfet$227
Xnfet$249_3 m1_n6433_17343# vss m1_n6274_17836# vss nfet$249
Xnfet$241_21 m1_28991_24224# m1_28991_24224# m1_28635_24542# m1_28635_24542# m1_29089_24542#
+ vss nfet$241
Xnfet$241_10 m1_17546_25658# m1_17546_25658# vss vss m1_18005_25502# vss nfet$241
Xnfet$247_0 m1_n3534_17714# vss m1_2384_19550# vss nfet$247
Xnfet$261_2 m1_9944_16080# m1_9944_16080# vss vss m1_11507_17358# vss nfet$261
Xnfet$254_1 m1_11671_21786# m1_11671_21786# vss vss m1_10509_21586# vss nfet$254
Xpfet$246_2 vdd m1_n4994_16080# m1_n5461_18030# m1_n6433_17343# pfet$246
Xpfet$253_3 vdd vdd m1_n4978_24224# vss pfet$253
Xpfet$239_1 vdd m1_n910_23922# m1_n646_24542# m1_n1271_25858# pfet$239
Xpfet$232_8 vdd vdd m1_28113_15778# m1_28470_16080# pfet$232
Xpfet$251_0 vdd vdd m1_n8625_26174# m1_n9336_24346# pfet$251
Xpfet$229_27 vdd m1_14422_22513# m1_14422_22513# m1_14022_22402# m1_14556_21786# m1_14556_21786#
+ pfet$229
Xpfet$229_16 vdd m1_24973_22513# m1_24973_22513# m1_23945_22102# m1_25739_21786# m1_25739_21786#
+ pfet$229
Xpfet$228_104 vdd vdd m1_14127_16080# m1_n7513_20152# pfet$228
Xpfet$230_5 vdd vdd vdd m1_n695_19850# m1_1103_20152# m1_1103_20152# pfet$230
Xpfet$231_17 vdd vdd m1_25739_21786# m1_25107_21786# pfet$231
Xnfet$244_10 m1_9015_17714# m1_9015_17714# vss vss m1_14005_20470# vss nfet$244
Xnfet$277_0 m1_n6839_20152# vss m1_n8145_21908# vss nfet$277
Xnfet$249_4 m1_n7247_17714# vss m1_n4377_15778# vss nfet$249
Xnfet$270_7 m1_n3541_23922# m1_n3541_23922# m1_n3651_26174# m1_n3651_26174# m1_n3415_25502#
+ vss nfet$270
Xnfet$241_22 m1_29607_24346# m1_29607_24346# vss vss m1_29089_24542# vss nfet$241
Xpfet$227_93 vdd m1_28991_24224# m1_30095_25658# m1_28010_25858# pfet$227
Xpfet$227_82 vdd vdd m1_21241_24346# m1_n7513_20152# pfet$227
Xpfet$227_71 vdd vdd m1_11039_21786# m1_11760_25858# pfet$227
Xpfet$227_60 vdd vdd m1_20126_25858# m1_21241_24346# pfet$227
Xnfet$241_11 m1_16442_24224# m1_16442_24224# m1_16086_24542# m1_16086_24542# m1_16540_24542#
+ vss nfet$241
Xnfet$247_1 m1_n3218_15478# vss m1_4620_20152# vss nfet$247
Xnfet$261_3 m1_11381_15778# m1_11381_15778# m1_11271_18030# m1_11271_18030# m1_11507_17358#
+ vss nfet$261
Xnfet$254_2 m1_8154_21786# m1_8154_21786# vss vss m1_6992_21586# vss nfet$254
Xpfet$246_3 vdd m1_n6172_16202# m1_n6657_17518# m1_n6274_17836# pfet$246
Xpfet$253_4 vdd vdd m1_n5571_25662# m1_n10452_25858# pfet$253
Xpfet$239_2 vdd m1_n290_24224# m1_814_25658# m1_n1271_25858# pfet$239
Xpfet$232_9 vdd vdd m1_29087_15778# m1_26217_17714# pfet$232
Xpfet$229_28 vdd m1_14422_22513# m1_14422_22513# m1_13394_22102# m1_15188_21786# m1_15188_21786#
+ pfet$229
Xpfet$229_17 vdd m1_21456_22513# m1_21456_22513# m1_21056_22402# m1_21590_21786# m1_21590_21786#
+ pfet$229
Xpfet$244_0 vdd m1_32818_20470# m1_32818_20470# m1_33050_19550# m1_30256_19792# m1_30256_19792#
+ pfet$244
Xnfet$247_10 m1_26063_15478# vss m1_29239_20152# vss nfet$247
Xpfet$251_1 vdd m1_n8625_26174# vdd m1_n8848_25658# pfet$251
Xpfet$228_105 vdd vdd m1_14258_17518# m1_13668_17714# pfet$228
Xpfet$230_6 vdd vdd vdd m1_6339_19850# m1_8137_20152# m1_8137_20152# pfet$230
Xnfet$244_11 m1_13198_17714# m1_13198_17714# vss vss m1_17522_20470# vss nfet$244
Xnfet$249_5 m1_n7247_17714# vss m1_n6657_17518# vss nfet$249
Xnfet$241_23 m1_25424_24346# m1_25424_24346# m1_24309_25858# m1_24309_25858# m1_26371_25502#
+ vss nfet$241
Xpfet$227_94 vdd m1_28492_25858# vdd m1_30095_25658# pfet$227
Xpfet$227_83 vdd m1_21729_25658# m1_22522_24542# m1_19781_25662# pfet$227
Xpfet$227_72 vdd m1_13363_25658# m1_14156_24542# m1_11415_25662# pfet$227
Xpfet$227_61 vdd m1_24452_24542# vdd m1_25424_24346# pfet$227
Xpfet$227_50 vdd vdd m1_20268_25662# m1_20126_25858# pfet$227
Xnfet$241_12 m1_17058_24346# m1_17058_24346# m1_15943_25858# m1_15943_25858# m1_18005_25502#
+ vss nfet$241
Xnfet$261_4 m1_10560_16202# m1_10560_16202# vss vss m1_10042_16398# vss nfet$261
Xpfet$246_4 vdd m1_28113_15778# m1_27292_16202# m1_27031_17343# pfet$246
Xpfet$239_3 vdd m1_814_25658# m1_1607_24542# m1_n1134_25662# pfet$239
Xnfet$247_2 m1_n7401_15478# vss m1_1103_20152# vss nfet$247
Xpfet$253_5 vdd vdd m1_n4847_25662# m1_n10452_25858# pfet$253
Xnfet$254_3 m1_7522_21786# m1_7522_21786# vss vss m1_6360_21586# vss nfet$254
Xnfet$252_0 pd1 vss m1_n1263_21786# vss nfet$252
Xpfet$237_0 vdd vdd vdd m1_33050_22344# m1_31535_22102# m1_31535_22102# pfet$237
Xnfet$247_11 m1_9331_15478# vss m1_15171_20152# vss nfet$247
Xpfet$244_1 vdd vdd vdd m1_33050_19550# m1_31535_19792# m1_31535_19792# pfet$244
Xpfet$251_2 vdd m1_n3651_26174# vdd m1_n4978_24224# pfet$251
Xpfet$229_29 vdd vdd vdd m1_14022_22402# m1_12805_21786# m1_12805_21786# pfet$229
Xpfet$229_18 vdd vdd vdd m1_24573_22402# m1_23356_21786# m1_23356_21786# pfet$229
Xpfet$228_106 vdd vdd m1_14482_17343# m1_17381_17714# pfet$228
Xpfet$230_7 vdd vdd vdd m1_6975_19550# m1_965_15478# m1_965_15478# pfet$230
Xnfet$244_12 m1_16452_19550# m1_16452_19550# vss vss m1_16890_20470# vss nfet$244
Xnfet$249_6 m1_n7247_17714# vss m1_n7383_17599# vss nfet$249
Xpfet$227_95 vdd vdd m1_28991_24224# m1_28371_23922# pfet$227
Xpfet$227_84 vdd vdd m1_23827_25858# m1_18073_21786# pfet$227
Xpfet$227_73 vdd m1_16086_24542# vdd m1_17058_24346# pfet$227
Xpfet$227_62 vdd vdd m1_24452_24542# m1_24808_24224# pfet$227
Xpfet$227_51 vdd vdd m1_20625_24224# m1_20005_23922# pfet$227
Xpfet$227_40 vdd vdd m1_11760_25858# m1_12875_24346# pfet$227
Xnfet$241_24 m1_30095_25658# m1_30095_25658# vss vss m1_30554_25502# vss nfet$241
Xnfet$241_13 m1_13363_25658# m1_13363_25658# vss vss m1_13822_25502# vss nfet$241
Xpfet$246_5 vdd m1_29087_15778# m1_28470_16080# m1_27190_17836# pfet$246
Xnfet$247_3 m1_649_17714# vss m1_5901_19550# vss nfet$247
Xnfet$261_5 m1_9944_16080# m1_9944_16080# m1_9485_17714# m1_9485_17714# m1_10042_16398#
+ vss nfet$261
Xpfet$253_6 vdd vdd m1_n4623_25487# fin pfet$253
Xnfet$254_4 m1_1120_21786# m1_1120_21786# vss vss m1_n42_21586# vss nfet$254
Xpfet$239_4 vdd m1_33174_24224# m1_34278_25658# m1_32193_25858# pfet$239
Xnfet$252_1 pd2 vss m1_2254_21786# vss nfet$252
Xnfet$245_0 m1_9485_17714# vss m1_9015_17714# vss nfet$245
Xpfet$244_2 vdd m1_32818_21586# m1_32818_21586# m1_33050_22344# m1_30256_22102# m1_30256_22102#
+ pfet$244
Xnfet$247_12 m1_13514_15478# vss m1_18688_20152# vss nfet$247
Xpfet$251_3 vdd vdd m1_n3651_26174# m1_n3541_23922# pfet$251
Xpfet$229_19 vdd m1_24973_22513# m1_24973_22513# m1_24573_22402# m1_25107_21786# m1_25107_21786#
+ pfet$229
Xpfet$228_107 vdd m1_15921_16080# m1_15454_18030# m1_14482_17343# pfet$228
Xpfet$230_8 vdd m1_9624_19404# m1_9624_19404# m1_10492_19550# m1_4832_17714# m1_4832_17714#
+ pfet$230
Xnfet$244_13 m1_19969_19550# m1_19969_19550# vss vss m1_20407_20470# vss nfet$244
Xnfet$269_10 vss vss m1_n4978_24224# vss nfet$269
Xnfet$249_7 m1_26217_17714# vss m1_26807_17518# vss nfet$249
Xpfet$227_96 vdd m1_28635_24542# vdd m1_29607_24346# pfet$227
Xpfet$227_85 vdd m1_24188_23922# m1_24452_24542# m1_23827_25858# pfet$227
Xpfet$227_74 vdd vdd m1_14556_21786# m1_15943_25858# pfet$227
Xpfet$227_63 vdd vdd m1_19781_25662# m1_19644_25858# pfet$227
Xpfet$227_52 vdd m1_20268_25662# m1_20005_23922# m1_19781_25662# pfet$227
Xpfet$227_41 vdd vdd m1_9288_21786# pd4 pfet$227
Xpfet$227_30 vdd vdd m1_2912_25858# m1_488_21786# pfet$227
Xnfet$275_0 m1_n927_19404# m1_n927_19404# vss vss m1_n6282_20470# vss nfet$275
Xnfet$241_25 m1_29607_24346# m1_29607_24346# m1_28492_25858# m1_28492_25858# m1_30554_25502#
+ vss nfet$241
Xnfet$241_14 m1_12875_24346# m1_12875_24346# m1_11760_25858# m1_11760_25858# m1_13822_25502#
+ vss nfet$241
Xnfet$247_4 m1_4832_17714# vss m1_9418_19550# vss nfet$247
Xnfet$261_6 m1_1578_16080# m1_1578_16080# vss vss m1_3141_17358# vss nfet$261
Xnfet$254_5 m1_4005_21786# m1_4005_21786# vss vss m1_2843_21586# vss nfet$254
Xpfet$239_5 vdd m1_32817_25662# m1_32554_23922# m1_32330_25662# pfet$239
Xpfet$246_6 vdd m1_28470_16080# m1_28003_18030# m1_27031_17343# pfet$246
Xpfet$253_7 vdd vdd m1_n3541_23922# m1_n3184_24224# pfet$253
Xnfet$252_2 pd9 vss m1_26873_21786# vss nfet$252
Xnfet$245_1 m1_9015_17714# vss m1_6116_17343# vss nfet$245
Xpfet$251_4 vdd m1_n10452_25858# vdd m1_n4362_24346# pfet$251
Xpfet$228_108 vdd vdd m1_15454_18030# m1_15564_15778# pfet$228
Xnfet$247_13 m1_13198_17714# vss m1_16452_19550# vss nfet$247
Xpfet$230_9 vdd m1_9624_19404# m1_9624_19404# m1_9856_19850# m1_9418_19550# m1_9418_19550#
+ pfet$230
Xpfet$242_0 vdd vdd vdd m1_36073_22344# define define pfet$242
Xnfet$244_14 m1_17381_17714# m1_17381_17714# vss vss m1_21039_20470# vss nfet$244
Xnfet$269_11 m1_n10452_25858# vss m1_n4847_25662# vss nfet$269
Xpfet$227_97 vdd vdd m1_21590_21786# m1_24309_25858# pfet$227
Xpfet$227_86 vdd m1_28634_25662# m1_28371_23922# m1_28147_25662# pfet$227
Xpfet$227_75 vdd vdd m1_19644_25858# m1_14556_21786# pfet$227
Xpfet$227_64 vdd vdd m1_22522_24542# m1_20126_25858# pfet$227
Xpfet$227_53 vdd m1_20625_24224# m1_21729_25658# m1_19644_25858# pfet$227
Xpfet$227_42 vdd m1_11760_25858# vdd m1_13363_25658# pfet$227
Xnfet$249_8 m1_n7513_20152# vss m1_26676_16080# vss nfet$249
Xpfet$227_31 vdd m1_3273_23922# m1_3537_24542# m1_2912_25858# pfet$227
Xpfet$227_20 vdd vdd m1_4509_24346# m1_n7513_20152# pfet$227
Xnfet$268_0 m1_n3822_20130# m1_n3822_20130# m1_n4485_20152# m1_n4485_20152# m1_n3724_20470#
+ vss nfet$268
Xnfet$275_1 m1_n2543_20130# m1_n2543_20130# m1_n5227_20152# m1_n5227_20152# m1_n2445_20470#
+ vss nfet$275
Xnfet$241_26 m1_25912_25658# m1_25912_25658# vss vss m1_26371_25502# vss nfet$241
Xnfet$241_15 m1_25424_24346# m1_25424_24346# vss vss m1_24906_24542# vss nfet$241
Xnfet$247_5 m1_965_15478# vss m1_8137_20152# vss nfet$247
Xnfet$261_7 m1_5761_16080# m1_5761_16080# m1_5302_17714# m1_5302_17714# m1_5859_16398#
+ vss nfet$261
Xnfet$254_6 m1_4637_21786# m1_4637_21786# vss vss m1_3475_21586# vss nfet$254
Xpfet$239_6 vdd m1_34278_25658# m1_35071_24542# m1_32330_25662# pfet$239
Xpfet$246_7 vdd m1_27292_16202# m1_26807_17518# m1_27190_17836# pfet$246
Xpfet$253_8 vdd vdd m1_n2567_23922# m1_n7320_25516# pfet$253
.ends

.subckt pfet$297 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$325 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$306 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$308 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt nfet$323 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt nfet$316 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$321 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$304 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$302 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt nfet$328 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$300 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$298 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$326 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt nfet$319 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$324 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$309 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$317 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$307 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt nfet$322 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$315 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$320 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt pfet$305 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt pfet$303 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$301 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$327 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt pfet$299 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$318 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_PFD_DFF_20250831$1 vss down up vdd fref fdiv
Xpfet$297_2 vdd m1_1095_n4045# m1_832_n5785# m1_n3885_n4045# pfet$297
Xnfet$325_2 m1_832_n8573# vss m1_1452_n8889# vss nfet$325
Xpfet$306_11 vdd vdd down m1_2779_n10883# pfet$306
Xpfet$297_3 vdd m1_2556_n4049# m1_3349_n5165# m1_n3885_n4045# pfet$297
Xnfet$325_3 vdd vss m1_1095_n11125# vss nfet$325
Xpfet$306_12 vdd m1_2556_n10129# m1_3349_n9089# m1_n3884_n11124# pfet$306
Xpfet$308_0 m1_n4677_n8889# vdd vdd m1_n1925_n10720# pfet$308
Xnfet$323_0 m1_n3885_n4045# vss m1_n3099_n4095# vss nfet$323
Xnfet$325_4 m1_n3884_n11124# m1_832_n8573# m1_1096_n9089# vss nfet$325
Xpfet$306_13 vdd vdd m1_n5427_n8573# m1_n4677_n8889# pfet$306
Xnfet$316_0 m1_2068_n5361# m1_2068_n5361# vss vss m1_1550_n5165# vss nfet$316
Xpfet$308_1 m1_n1925_n10720# vdd vdd m1_n3098_n10720# pfet$308
Xnfet$323_1 m1_n3885_n6084# vss m1_n3099_n5680# vss nfet$323
Xnfet$325_5 m1_2758_n8889# vss m1_2068_n8889# vss nfet$325
Xpfet$306_14 vdd vdd m1_n3884_n11124# m1_n5427_n10882# pfet$306
Xnfet$316_1 m1_1452_n5483# m1_1452_n5483# m1_1096_n5165# m1_1096_n5165# m1_1550_n5165#
+ vss nfet$316
Xpfet$308_2 m1_n4677_n10522# vdd vdd m1_n1925_n9135# pfet$308
Xpfet$306_15 vdd m1_n5427_n10882# vdd m1_n5649_n11124# pfet$306
Xnfet$316_2 m1_2556_n4049# m1_2556_n4049# vss vss m1_3015_n4205# vss nfet$316
Xnfet$325_6 m1_2779_n10883# vss down vss nfet$325
Xpfet$308_3 m1_n1925_n9135# vdd vdd m1_n3098_n9135# pfet$308
Xpfet$306_0 vdd vdd m1_2779_n10883# m1_2068_n8889# pfet$306
Xnfet$321_0 m1_n5428_n3533# vss m1_n3885_n4045# vss nfet$321
Xnfet$325_7 m1_2779_n10883# vss m1_3349_n9089# vss nfet$325
Xpfet$306_16 vdd vdd m1_n5427_n10882# m1_n4677_n10522# pfet$306
Xnfet$316_3 m1_2068_n5361# m1_2068_n5361# m1_2779_n3533# m1_2779_n3533# m1_3015_n4205#
+ vss nfet$316
Xnfet$321_1 m1_n5868_n3849# vss m1_n5650_n4045# vss nfet$321
Xpfet$306_1 vdd m1_2779_n10883# vdd m1_2556_n10129# pfet$306
Xpfet$306_17 vdd vdd m1_n5649_n11124# m1_n5867_n10544# pfet$306
Xnfet$325_8 m1_n3884_n9085# m1_2556_n10129# m1_3349_n9089# vss nfet$325
Xpfet$306_2 vdd m1_1095_n11125# m1_832_n8573# m1_n3884_n11124# pfet$306
Xnfet$321_2 m1_n5428_n5842# vss m1_n3885_n6084# vss nfet$321
Xnfet$325_9 m1_n5427_n10882# vss m1_n3884_n11124# vss nfet$325
Xpfet$306_18 vdd vdd m1_n5867_n10544# fdiv pfet$306
Xpfet$306_3 vdd m1_1452_n8889# m1_2556_n10129# m1_n3884_n9085# pfet$306
Xpfet$304_0 vdd m1_n5428_n3533# vdd m1_n5650_n4045# pfet$304
Xnfet$321_3 fref vss m1_n5868_n3849# vss nfet$321
Xpfet$306_19 vdd vdd m1_n3884_n9085# m1_n5427_n8573# pfet$306
Xpfet$306_4 vdd vdd m1_1452_n8889# m1_832_n8573# pfet$306
Xpfet$304_1 vdd vdd m1_n5428_n3533# m1_n4678_n3849# pfet$304
Xpfet$306_5 vdd vdd m1_1095_n11125# vdd pfet$306
Xpfet$304_2 vdd m1_n5428_n5842# vdd m1_n5868_n3849# pfet$304
Xpfet$306_6 vdd vdd m1_1096_n9089# m1_1452_n8889# pfet$306
Xpfet$304_3 vdd vdd m1_n5428_n5842# m1_n4678_n5482# pfet$304
Xpfet$302_0 m1_n1926_n4095# vdd vdd m1_n3099_n4095# pfet$302
Xnfet$328_0 up up m1_5895_n8089# m1_5895_n8089# m1_5043_n9245# vss nfet$328
Xpfet$306_7 vdd m1_832_n8573# m1_1096_n9089# m1_n3884_n9085# pfet$306
Xpfet$302_1 m1_n4678_n3849# vdd vdd m1_n1926_n5680# pfet$302
Xnfet$328_1 down down vss vss m1_5043_n9245# vss nfet$328
Xpfet$306_8 vdd m1_1096_n9089# vdd m1_2068_n8889# pfet$306
Xpfet$302_2 m1_n1926_n5680# vdd vdd m1_n3099_n5680# pfet$302
Xpfet$306_9 vdd vdd m1_2068_n8889# m1_2758_n8889# pfet$306
Xpfet$302_3 m1_n4678_n5482# vdd vdd m1_n1926_n4095# pfet$302
Xpfet$300_0 vdd vdd m1_2758_n8889# m1_4978_n5483# pfet$300
Xpfet$298_0 vdd vdd m1_1096_n5165# m1_1452_n5483# pfet$298
Xnfet$326_0 m1_n3884_n11124# vss m1_n3098_n10720# vss nfet$326
Xpfet$298_1 vdd m1_1096_n5165# vdd m1_2068_n5361# pfet$298
Xnfet$326_1 m1_n3884_n9085# vss m1_n3098_n9135# vss nfet$326
Xnfet$319_0 m1_5895_n8089# vss m1_5464_n5483# vss nfet$319
Xpfet$298_2 vdd m1_2779_n3533# vdd m1_2556_n4049# pfet$298
Xnfet$319_1 m1_5464_n5483# vss m1_4978_n5483# vss nfet$319
Xpfet$298_3 vdd vdd m1_2779_n3533# m1_2068_n5361# pfet$298
Xnfet$324_0 m1_2556_n10129# m1_2556_n10129# vss vss m1_3015_n10205# vss nfet$324
Xpfet$309_0 vdd m1_5895_n8089# vdd down pfet$309
Xnfet$325_10 m1_n5867_n10544# vss m1_n5649_n11124# vss nfet$325
Xnfet$324_1 m1_1452_n8889# m1_1452_n8889# m1_1096_n9089# m1_1096_n9089# m1_1550_n9245#
+ vss nfet$324
Xpfet$309_1 vdd vdd m1_5895_n8089# up pfet$309
Xnfet$317_0 m1_2779_n3533# vss up vss nfet$317
Xnfet$325_11 fdiv vss m1_n5867_n10544# vss nfet$325
Xnfet$324_2 m1_2068_n8889# m1_2068_n8889# vss vss m1_1550_n9245# vss nfet$324
Xnfet$317_1 m1_2779_n3533# vss m1_3349_n5165# vss nfet$317
Xnfet$325_12 m1_n5427_n8573# vss m1_n3884_n9085# vss nfet$325
Xnfet$317_2 m1_2758_n8889# vss m1_2068_n5361# vss nfet$317
Xnfet$324_3 m1_2068_n8889# m1_2068_n8889# m1_2779_n10883# m1_2779_n10883# m1_3015_n10205#
+ vss nfet$324
Xpfet$307_0 vdd vdd m1_n3098_n10720# m1_n3884_n11124# pfet$307
Xnfet$322_0 m1_n4678_n3849# m1_n4678_n3849# m1_n5428_n3533# m1_n5428_n3533# m1_n5192_n4205#
+ vss nfet$322
Xnfet$317_3 m1_832_n5785# vss m1_1452_n5483# vss nfet$317
Xnfet$324_4 m1_n4677_n10522# m1_n4677_n10522# m1_n5427_n10882# m1_n5427_n10882# m1_n5191_n10204#
+ vss nfet$324
Xnfet$315_0 m1_n3885_n4045# m1_832_n5785# m1_1096_n5165# vss nfet$315
Xpfet$307_1 vdd vdd m1_n3098_n9135# m1_n3884_n9085# pfet$307
Xnfet$322_1 m1_n5650_n4045# m1_n5650_n4045# vss vss m1_n5192_n4205# vss nfet$322
Xnfet$317_4 vdd vss m1_1095_n4045# vss nfet$317
Xnfet$315_1 m1_n3885_n4045# m1_1452_n5483# m1_2556_n4049# vss nfet$315
Xnfet$324_5 m1_n5649_n11124# m1_n5649_n11124# vss vss m1_n5191_n10204# vss nfet$324
Xnfet$322_2 m1_n4678_n5482# m1_n4678_n5482# m1_n5428_n5842# m1_n5428_n5842# m1_n5192_n5164#
+ vss nfet$322
Xnfet$324_6 m1_n4677_n8889# m1_n4677_n8889# m1_n5427_n8573# m1_n5427_n8573# m1_n5191_n9245#
+ vss nfet$324
Xnfet$315_2 m1_n3885_n6084# m1_1095_n4045# m1_832_n5785# vss nfet$315
Xnfet$322_3 m1_n5868_n3849# m1_n5868_n3849# vss vss m1_n5192_n5164# vss nfet$322
Xnfet$320_0 m1_n1926_n4095# m1_n3099_n4095# vss vss nfet$320
Xpfet$305_0 vdd vdd m1_n3099_n4095# m1_n3885_n4045# pfet$305
Xnfet$315_3 m1_n3885_n6084# m1_2556_n4049# m1_3349_n5165# vss nfet$315
Xnfet$324_7 m1_n5867_n10544# m1_n5867_n10544# vss vss m1_n5191_n9245# vss nfet$324
Xnfet$320_1 m1_n4678_n3849# m1_n1926_n5680# vss vss nfet$320
Xpfet$305_1 vdd vdd m1_n3099_n5680# m1_n3885_n6084# pfet$305
Xnfet$320_2 m1_n1926_n5680# m1_n3099_n5680# vss vss nfet$320
Xnfet$320_3 m1_n4678_n5482# m1_n1926_n4095# vss vss nfet$320
Xpfet$303_0 vdd vdd m1_n3885_n4045# m1_n5428_n3533# pfet$303
Xpfet$303_1 vdd vdd m1_n5650_n4045# m1_n5868_n3849# pfet$303
Xpfet$303_2 vdd vdd m1_n3885_n6084# m1_n5428_n5842# pfet$303
Xpfet$303_3 vdd vdd m1_n5868_n3849# fref pfet$303
Xpfet$301_0 vdd vdd m1_5464_n5483# m1_5895_n8089# pfet$301
Xnfet$327_0 m1_n4677_n8889# m1_n1925_n10720# vss vss nfet$327
Xpfet$299_0 vdd vdd m1_3349_n5165# m1_2779_n3533# pfet$299
Xpfet$301_1 vdd vdd m1_4978_n5483# m1_5464_n5483# pfet$301
Xpfet$299_1 vdd vdd up m1_2779_n3533# pfet$299
Xnfet$327_1 m1_n1925_n10720# m1_n3098_n10720# vss vss nfet$327
Xpfet$299_2 vdd vdd m1_2068_n5361# m1_2758_n8889# pfet$299
Xnfet$327_2 m1_n4677_n10522# m1_n1925_n9135# vss vss nfet$327
Xpfet$299_3 vdd vdd m1_1452_n5483# m1_832_n5785# pfet$299
Xpfet$297_0 vdd m1_832_n5785# m1_1096_n5165# m1_n3885_n6084# pfet$297
Xnfet$325_0 m1_n3884_n9085# m1_1095_n11125# m1_832_n8573# vss nfet$325
Xnfet$327_3 m1_n1925_n9135# m1_n3098_n9135# vss vss nfet$327
Xpfet$306_20 vdd m1_n5427_n8573# vdd m1_n5867_n10544# pfet$306
Xpfet$299_4 vdd vdd m1_1095_n4045# vdd pfet$299
Xpfet$297_1 vdd m1_1452_n5483# m1_2556_n4049# m1_n3885_n6084# pfet$297
Xnfet$325_1 m1_n3884_n11124# m1_1452_n8889# m1_2556_n10129# vss nfet$325
Xpfet$306_10 vdd vdd m1_3349_n9089# m1_2779_n10883# pfet$306
Xnfet$318_0 m1_4978_n5483# vss m1_2758_n8889# vss nfet$318
.ends

.subckt asc_drive_buffer$2 vss in vdd out
Xpfet$295_0 vdd vdd m1_4002_n1060# m1_3466_n454# pfet$295
Xpfet$293_0 out out m1_4274_n1060# vdd m1_4274_n1060# out vdd vdd m1_4274_n1060# out
+ m1_4274_n1060# m1_4274_n1060# out m1_4274_n1060# vdd m1_4274_n1060# vdd m1_4274_n1060#
+ pfet$293
Xnfet$314_0 in vss m1_3466_n454# vss nfet$314
Xnfet$312_0 out out vss m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# m1_4274_n1060#
+ m1_4274_n1060# out m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# vss vss
+ nfet$312
Xpfet$296_0 vdd vdd m1_3466_n454# in pfet$296
Xpfet$294_0 m1_4274_n1060# vdd vdd m1_4274_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ vdd m1_4002_n1060# m1_4002_n1060# pfet$294
Xnfet$313_0 m1_3466_n454# vss m1_4002_n1060# vss nfet$313
Xnfet$311_0 m1_4274_n1060# vss m1_4002_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ m1_4274_n1060# vss m1_4002_n1060# vss nfet$311
.ends

.subckt pfet$288 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$309 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$307 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$291 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$310 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$289 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$308 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$292 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$306 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$290 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt asc_drive_buffer_up$1 vss out in vdd
Xpfet$288_0 out out m1_778_712# vdd m1_778_712# out vdd vdd m1_778_712# out m1_778_712#
+ m1_778_712# out m1_778_712# vdd m1_778_712# vdd m1_778_712# pfet$288
Xnfet$309_0 m1_n566_1318# vss m1_n30_1318# vss nfet$309
Xnfet$307_0 out out vss m1_778_712# m1_778_712# out vss m1_778_712# m1_778_712# m1_778_712#
+ out m1_778_712# m1_778_712# out vss m1_778_712# vss vss nfet$307
Xpfet$291_0 vdd vdd m1_n30_1318# m1_n566_1318# pfet$291
Xnfet$310_0 in vss m1_n566_1318# vss nfet$310
Xpfet$289_0 m1_778_712# vdd vdd m1_778_712# m1_506_712# m1_506_712# m1_778_712# vdd
+ m1_506_712# m1_506_712# pfet$289
Xnfet$308_0 m1_n30_1318# vss m1_506_712# vss nfet$308
Xpfet$292_0 vdd vdd m1_n566_1318# in pfet$292
Xnfet$306_0 m1_778_712# vss m1_506_712# m1_506_712# m1_506_712# m1_778_712# m1_778_712#
+ vss m1_506_712# vss nfet$306
Xpfet$290_0 vdd vdd m1_506_712# m1_n30_1318# pfet$290
.ends

.subckt pfet$310 a_254_0# a_348_560# w_n180_n88# a_414_0# a_n92_0# a_94_0# a_574_0#
+ a_508_560# a_188_560# a_28_560#
X0 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$329 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt BIAS$1 vdd vss 100n 200n res 200p1 200p2
Xpfet$310_10 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$310
Xpfet$310_11 vdd res vdd 200n vdd 200n vdd res res res pfet$310
Xpfet$310_12 vdd res vdd 100n vdd 100n vdd res res res pfet$310
Xpfet$310_13 vdd res vdd res vdd res vdd res res res pfet$310
Xpfet$310_0 vdd res vdd 200n vdd 200n vdd res res res pfet$310
Xpfet$310_15 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$310
Xpfet$310_14 vdd res vdd 200n vdd 200n vdd res res res pfet$310
Xpfet$310_1 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$310
Xpfet$310_2 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$310
Xnfet$329_1 vss vss vss vss vss vss vss vss vss vss nfet$329
Xnfet$329_0 m1_27_n1423# vss 200p1 m1_27_n1423# vss 200p1 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$329
Xpfet$310_3 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$310
Xnfet$329_2 m1_27_n1423# vss 200p2 m1_27_n1423# vss 200p2 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$329
Xpfet$310_4 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$310
Xnfet$329_3 vss vss vss vss vss vss vss vss vss vss nfet$329
Xpfet$310_5 vdd res vdd 200n vdd 200n vdd res res res pfet$310
Xnfet$329_4 m1_27_n1423# vss 200p2 m1_27_n1423# vss 200p2 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$329
Xpfet$310_7 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$310
Xpfet$310_6 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$310
Xnfet$329_5 m1_27_n1423# vss 200p1 m1_27_n1423# vss 200p1 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$329
Xnfet$329_6 m1_27_n1423# vss m1_27_n1423# m1_27_n1423# vss m1_27_n1423# m1_27_n1423#
+ vss m1_27_n1423# vss nfet$329
Xpfet$310_8 vdd res vdd res vdd res vdd res res res pfet$310
Xnfet$329_7 m1_27_n1423# vss m1_27_n1423# m1_27_n1423# vss m1_27_n1423# m1_27_n1423#
+ vss m1_27_n1423# vss nfet$329
Xpfet$310_9 vdd res vdd 100n vdd 100n vdd res res res pfet$310
.ends

.subckt nfet$300 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$291 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$276 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$298 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$274 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$272 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$296 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$289 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$294 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$279 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$284 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$292 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$277 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$282 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$275 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$290 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt nfet$303 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$280 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$273 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$301 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$299 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$271 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$297 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$295 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$285 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$293 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$278 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$283 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$281 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$302 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_lock_detector_20250826$1 ref vdd div lock vss
Xnfet$300_0 div m1_n4030_5270# vss vss nfet$300
Xnfet$291_7 m1_3254_4493# vss m1_2982_4493# m1_2982_4493# m1_2982_4493# m1_3254_4493#
+ m1_3254_4493# vss m1_2982_4493# vss nfet$291
Xpfet$276_7 vdd m1_16242_6960# m1_15979_5220# m1_15755_6960# pfet$276
Xnfet$298_0 m1_15979_2344# vss m1_16599_2028# vss nfet$298
Xpfet$274_4 m1_n940_4493# vdd vdd m1_n940_4493# m1_n1212_4493# m1_n1212_4493# m1_n940_4493#
+ vdd m1_n1212_4493# m1_n1212_4493# pfet$274
Xpfet$272_1 vdd vdd m1_11370_n340# m1_10834_1478# pfet$272
Xnfet$300_1 m1_n6066_7868# vss m1_n4030_5270# vss nfet$300
Xnfet$298_1 m1_15618_394# vss m1_15755_n208# vss nfet$298
Xpfet$274_5 m1_11642_4493# vdd vdd m1_11642_4493# m1_11370_4493# m1_11370_4493# m1_11642_4493#
+ vdd m1_11370_4493# m1_11370_4493# pfet$274
Xpfet$272_2 vdd vdd m1_2982_n340# m1_2446_1478# pfet$272
Xnfet$298_2 m1_n2336_5099# vss m1_16242_n208# vss nfet$298
Xpfet$274_6 m1_3254_4493# vdd vdd m1_3254_4493# m1_2982_4493# m1_2982_4493# m1_3254_4493#
+ vdd m1_2982_4493# m1_2982_4493# pfet$274
Xpfet$272_3 vdd vdd m1_n1212_n340# m1_n1748_1478# pfet$272
Xnfet$298_3 m1_17926_34# vss m1_18496_1828# vss nfet$298
Xnfet$296_0 m1_15755_n208# m1_16599_2028# m1_17703_788# vss nfet$296
Xpfet$274_7 m1_7448_4493# vdd vdd m1_7448_4493# m1_7176_4493# m1_7176_4493# m1_7448_4493#
+ vdd m1_7176_4493# m1_7176_4493# pfet$274
Xpfet$272_4 vdd vdd m1_n1212_4493# m1_n1748_5099# pfet$272
Xnfet$298_4 m1_12790_n340# vss m1_15618_394# vss nfet$298
Xnfet$296_1 m1_15618_394# m1_16242_n208# m1_15979_2344# vss nfet$296
Xnfet$289_0 m1_8596_n340# m1_8596_n340# vss m1_7448_n340# m1_7448_n340# m1_8596_n340#
+ vss m1_7448_n340# m1_7448_n340# m1_7448_n340# m1_8596_n340# m1_7448_n340# m1_7448_n340#
+ m1_8596_n340# vss m1_7448_n340# vss vss nfet$289
Xpfet$272_5 vdd vdd m1_2982_4493# m1_2446_5099# pfet$272
Xnfet$289_1 m1_4402_n340# m1_4402_n340# vss m1_3254_n340# m1_3254_n340# m1_4402_n340#
+ vss m1_3254_n340# m1_3254_n340# m1_3254_n340# m1_4402_n340# m1_3254_n340# m1_3254_n340#
+ m1_4402_n340# vss m1_3254_n340# vss vss nfet$289
Xnfet$296_2 m1_15618_394# m1_17703_788# m1_18496_1828# vss nfet$296
Xnfet$298_5 vss vss m1_17215_2028# vss nfet$298
Xpfet$272_6 vdd vdd m1_7176_4493# m1_6640_5099# pfet$272
Xnfet$298_6 m1_17926_34# vss m1_19469_1832# vss nfet$298
Xnfet$294_0 m1_n7214_4493# vss m1_n7486_4493# m1_n7486_4493# m1_n7486_4493# m1_n7214_4493#
+ m1_n7214_4493# vss m1_n7486_4493# vss nfet$294
Xnfet$289_2 m1_12790_n340# m1_12790_n340# vss m1_11642_n340# m1_11642_n340# m1_12790_n340#
+ vss m1_11642_n340# m1_11642_n340# m1_11642_n340# m1_12790_n340# m1_11642_n340# m1_11642_n340#
+ m1_12790_n340# vss m1_11642_n340# vss vss nfet$289
Xnfet$296_3 m1_15755_n208# m1_15979_2344# m1_16243_1828# vss nfet$296
Xpfet$272_7 vdd vdd m1_11370_4493# m1_10834_5099# pfet$272
Xpfet$279_0 m1_n11408_4493# vdd vdd m1_n11408_4493# m1_n11680_4493# m1_n11680_4493#
+ m1_n11408_4493# vdd m1_n11680_4493# m1_n11680_4493# pfet$279
Xnfet$296_4 m1_15618_7156# m1_17703_6956# m1_18496_5840# vss nfet$296
Xnfet$289_3 m1_208_n340# m1_208_n340# vss m1_n940_n340# m1_n940_n340# m1_208_n340#
+ vss m1_n940_n340# m1_n940_n340# m1_n940_n340# m1_208_n340# m1_n940_n340# m1_n940_n340#
+ m1_208_n340# vss m1_n940_n340# vss vss nfet$289
Xnfet$298_7 vss vss m1_17215_5644# vss nfet$298
Xnfet$294_1 m1_n15602_4493# vss m1_n15874_4493# m1_n15874_4493# m1_n15874_4493# m1_n15602_4493#
+ m1_n15602_4493# vss m1_n15874_4493# vss nfet$294
Xpfet$279_1 m1_n7214_4493# vdd vdd m1_n7214_4493# m1_n7486_4493# m1_n7486_4493# m1_n7214_4493#
+ vdd m1_n7486_4493# m1_n7486_4493# pfet$279
Xnfet$298_8 m1_17926_7472# vss m1_19469_4920# vss nfet$298
Xnfet$289_4 m1_12790_7868# m1_12790_7868# vss m1_11642_4493# m1_11642_4493# m1_12790_7868#
+ vss m1_11642_4493# m1_11642_4493# m1_11642_4493# m1_12790_7868# m1_11642_4493# m1_11642_4493#
+ m1_12790_7868# vss m1_11642_4493# vss vss nfet$289
Xnfet$296_5 m1_15755_6960# m1_15979_5220# m1_16243_5840# vss nfet$296
Xnfet$294_2 m1_n11408_4493# vss m1_n11680_4493# m1_n11680_4493# m1_n11680_4493# m1_n11408_4493#
+ m1_n11408_4493# vss m1_n11680_4493# vss nfet$294
Xpfet$284_0 vdd m1_19675_2344# vdd m1_19469_1832# pfet$284
Xpfet$279_2 m1_n15602_4493# vdd vdd m1_n15602_4493# m1_n15874_4493# m1_n15874_4493#
+ m1_n15602_4493# vdd m1_n15874_4493# m1_n15874_4493# pfet$279
Xnfet$289_5 m1_8596_7868# m1_8596_7868# vss m1_7448_4493# m1_7448_4493# m1_8596_7868#
+ vss m1_7448_4493# m1_7448_4493# m1_7448_4493# m1_8596_7868# m1_7448_4493# m1_7448_4493#
+ m1_8596_7868# vss m1_7448_4493# vss vss nfet$289
Xnfet$296_6 m1_15618_7156# m1_16242_6960# m1_15979_5220# vss nfet$296
Xnfet$298_9 m1_17926_7472# vss m1_18496_5840# vss nfet$298
Xnfet$292_0 m1_n6066_7868# m1_n6066_7868# vss m1_n7214_4493# m1_n7214_4493# m1_n6066_7868#
+ vss m1_n7214_4493# m1_n7214_4493# m1_n7214_4493# m1_n6066_7868# m1_n7214_4493# m1_n7214_4493#
+ m1_n6066_7868# vss m1_n7214_4493# vss vss nfet$292
Xpfet$277_0 vdd m1_17926_34# vdd m1_17703_788# pfet$277
Xpfet$284_1 vdd vdd m1_19675_2344# m1_19469_4920# pfet$284
Xnfet$289_6 m1_208_7868# m1_208_7868# vss m1_n940_4493# m1_n940_4493# m1_208_7868#
+ vss m1_n940_4493# m1_n940_4493# m1_n940_4493# m1_208_7868# m1_n940_4493# m1_n940_4493#
+ m1_208_7868# vss m1_n940_4493# vss vss nfet$289
Xnfet$296_7 m1_15755_6960# m1_16599_5522# m1_17703_6956# vss nfet$296
Xnfet$292_1 m1_n14454_7868# m1_n14454_7868# vss m1_n15602_4493# m1_n15602_4493# m1_n14454_7868#
+ vss m1_n15602_4493# m1_n15602_4493# m1_n15602_4493# m1_n14454_7868# m1_n15602_4493#
+ m1_n15602_4493# m1_n14454_7868# vss m1_n15602_4493# vss vss nfet$292
Xpfet$277_1 vdd vdd m1_17926_34# m1_17215_2028# pfet$277
Xnfet$289_7 m1_4402_7868# m1_4402_7868# vss m1_3254_4493# m1_3254_4493# m1_4402_7868#
+ vss m1_3254_4493# m1_3254_4493# m1_3254_4493# m1_4402_7868# m1_3254_4493# m1_3254_4493#
+ m1_4402_7868# vss m1_3254_4493# vss vss nfet$289
Xnfet$292_2 m1_n10260_7868# m1_n10260_7868# vss m1_n11408_4493# m1_n11408_4493# m1_n10260_7868#
+ vss m1_n11408_4493# m1_n11408_4493# m1_n11408_4493# m1_n10260_7868# m1_n11408_4493#
+ m1_n11408_4493# m1_n10260_7868# vss m1_n11408_4493# vss vss nfet$292
Xpfet$277_2 vdd m1_16243_1828# vdd m1_17215_2028# pfet$277
Xpfet$282_0 vdd vdd vdd m1_n3798_6028# div div pfet$282
Xpfet$275_0 vdd vdd m1_16599_2028# m1_15979_2344# pfet$275
Xnfet$290_0 m1_10834_1478# vss m1_11370_n340# vss nfet$290
Xpfet$277_3 vdd vdd m1_16243_1828# m1_16599_2028# pfet$277
Xpfet$282_1 vdd m1_n4030_5270# m1_n4030_5270# m1_n3798_6028# m1_n6066_7868# m1_n6066_7868#
+ pfet$282
Xnfet$303_0 m1_19675_2344# vss lock vss nfet$303
Xpfet$277_4 vdd m1_16243_5840# vdd m1_17215_5644# pfet$277
Xpfet$275_1 vdd vdd m1_16242_n208# m1_n2336_5099# pfet$275
Xnfet$290_1 m1_2446_1478# vss m1_2982_n340# vss nfet$290
Xpfet$277_5 vdd vdd m1_16243_5840# m1_16599_5522# pfet$277
Xpfet$275_2 vdd vdd m1_15755_n208# m1_15618_394# pfet$275
Xnfet$290_2 m1_6640_1478# vss m1_7176_n340# vss nfet$290
Xpfet$280_0 vdd vdd m1_n11680_4493# m1_n12216_5099# pfet$280
Xpfet$277_6 vdd m1_17926_7472# vdd m1_17703_6956# pfet$277
Xpfet$275_3 vdd vdd m1_18496_1828# m1_17926_34# pfet$275
Xnfet$290_3 m1_n1748_1478# vss m1_n1212_n340# vss nfet$290
Xpfet$273_0 m1_8596_n340# m1_8596_n340# m1_7448_n340# vdd m1_7448_n340# m1_8596_n340#
+ vdd vdd m1_7448_n340# m1_8596_n340# m1_7448_n340# m1_7448_n340# m1_8596_n340# m1_7448_n340#
+ vdd m1_7448_n340# vdd m1_7448_n340# pfet$273
Xnfet$301_0 m1_n4030_5270# vss m1_n2336_5099# vss nfet$301
Xpfet$280_1 vdd vdd m1_n7486_4493# m1_n8022_5099# pfet$280
Xnfet$299_0 m1_n14454_7868# vss m1_n12216_5099# vss nfet$299
Xnfet$290_4 m1_10834_5099# vss m1_11370_4493# vss nfet$290
Xpfet$277_7 vdd vdd m1_17926_7472# m1_17215_5644# pfet$277
Xpfet$275_4 vdd vdd m1_15618_394# m1_12790_n340# pfet$275
Xpfet$273_1 m1_12790_n340# m1_12790_n340# m1_11642_n340# vdd m1_11642_n340# m1_12790_n340#
+ vdd vdd m1_11642_n340# m1_12790_n340# m1_11642_n340# m1_11642_n340# m1_12790_n340#
+ m1_11642_n340# vdd m1_11642_n340# vdd m1_11642_n340# pfet$273
Xpfet$280_2 vdd vdd m1_n15874_4493# m1_n16410_5099# pfet$280
Xnfet$299_1 div vss m1_n16410_5099# vss nfet$299
Xnfet$290_5 m1_6640_5099# vss m1_7176_4493# vss nfet$290
Xpfet$275_5 vdd vdd m1_17215_2028# vss pfet$275
Xpfet$273_2 m1_4402_n340# m1_4402_n340# m1_3254_n340# vdd m1_3254_n340# m1_4402_n340#
+ vdd vdd m1_3254_n340# m1_4402_n340# m1_3254_n340# m1_3254_n340# m1_4402_n340# m1_3254_n340#
+ vdd m1_3254_n340# vdd m1_3254_n340# pfet$273
Xnfet$299_2 m1_n10260_7868# vss m1_n8022_5099# vss nfet$299
Xnfet$290_6 m1_n1748_5099# vss m1_n1212_4493# vss nfet$290
Xpfet$275_6 vdd vdd m1_19469_1832# m1_17926_34# pfet$275
Xpfet$273_3 m1_208_n340# m1_208_n340# m1_n940_n340# vdd m1_n940_n340# m1_208_n340#
+ vdd vdd m1_n940_n340# m1_208_n340# m1_n940_n340# m1_n940_n340# m1_208_n340# m1_n940_n340#
+ vdd m1_n940_n340# vdd m1_n940_n340# pfet$273
Xpfet$271_0 vdd vdd m1_6640_1478# m1_4402_n340# pfet$271
Xnfet$297_0 m1_17215_2028# m1_17215_2028# m1_17926_34# m1_17926_34# m1_18162_712#
+ vss nfet$297
Xnfet$290_7 m1_2446_5099# vss m1_2982_4493# vss nfet$290
Xpfet$275_7 vdd vdd m1_17215_5644# vss pfet$275
Xpfet$271_1 vdd vdd m1_10834_1478# m1_8596_n340# pfet$271
Xpfet$273_4 m1_208_7868# m1_208_7868# m1_n940_4493# vdd m1_n940_4493# m1_208_7868#
+ vdd vdd m1_n940_4493# m1_208_7868# m1_n940_4493# m1_n940_4493# m1_208_7868# m1_n940_4493#
+ vdd m1_n940_4493# vdd m1_n940_4493# pfet$273
Xnfet$297_1 m1_17703_788# m1_17703_788# vss vss m1_18162_712# vss nfet$297
Xpfet$273_5 m1_12790_7868# m1_12790_7868# m1_11642_4493# vdd m1_11642_4493# m1_12790_7868#
+ vdd vdd m1_11642_4493# m1_12790_7868# m1_11642_4493# m1_11642_4493# m1_12790_7868#
+ m1_11642_4493# vdd m1_11642_4493# vdd m1_11642_4493# pfet$273
Xpfet$275_8 vdd vdd m1_19469_4920# m1_17926_7472# pfet$275
Xpfet$271_2 vdd vdd m1_n1748_1478# ref pfet$271
Xpfet$275_9 vdd vdd m1_18496_5840# m1_17926_7472# pfet$275
Xnfet$297_2 m1_16599_2028# m1_16599_2028# m1_16243_1828# m1_16243_1828# m1_16697_1672#
+ vss nfet$297
Xpfet$273_6 m1_4402_7868# m1_4402_7868# m1_3254_4493# vdd m1_3254_4493# m1_4402_7868#
+ vdd vdd m1_3254_4493# m1_4402_7868# m1_3254_4493# m1_3254_4493# m1_4402_7868# m1_3254_4493#
+ vdd m1_3254_4493# vdd m1_3254_4493# pfet$273
Xpfet$271_3 vdd vdd m1_n1748_5099# m1_n2336_5099# pfet$271
Xnfet$297_3 m1_17215_2028# m1_17215_2028# vss vss m1_16697_1672# vss nfet$297
Xpfet$273_7 m1_8596_7868# m1_8596_7868# m1_7448_4493# vdd m1_7448_4493# m1_8596_7868#
+ vdd vdd m1_7448_4493# m1_8596_7868# m1_7448_4493# m1_7448_4493# m1_8596_7868# m1_7448_4493#
+ vdd m1_7448_4493# vdd m1_7448_4493# pfet$273
Xnfet$295_0 m1_8596_n340# vss m1_10834_1478# vss nfet$295
Xpfet$271_4 vdd vdd m1_6640_5099# m1_4402_7868# pfet$271
Xnfet$295_1 m1_4402_n340# vss m1_6640_1478# vss nfet$295
Xnfet$297_4 m1_17215_5644# m1_17215_5644# vss vss m1_16697_5840# vss nfet$297
Xpfet$271_5 vdd vdd m1_10834_5099# m1_8596_7868# pfet$271
Xnfet$297_5 m1_16599_5522# m1_16599_5522# m1_16243_5840# m1_16243_5840# m1_16697_5840#
+ vss nfet$297
Xnfet$298_10 m1_12790_7868# vss m1_15618_7156# vss nfet$298
Xnfet$295_2 ref vss m1_n1748_1478# vss nfet$295
Xpfet$271_6 vdd vdd m1_2446_5099# m1_208_7868# pfet$271
Xpfet$285_0 vdd vdd lock m1_19675_2344# pfet$285
Xnfet$297_6 m1_17215_5644# m1_17215_5644# m1_17926_7472# m1_17926_7472# m1_18162_6800#
+ vss nfet$297
Xnfet$298_11 m1_15979_5220# vss m1_16599_5522# vss nfet$298
Xnfet$295_3 m1_n2336_5099# vss m1_n1748_5099# vss nfet$295
Xnfet$293_0 m1_n8022_5099# vss m1_n7486_4493# vss nfet$293
Xpfet$278_0 m1_n10260_7868# m1_n10260_7868# m1_n11408_4493# vdd m1_n11408_4493# m1_n10260_7868#
+ vdd vdd m1_n11408_4493# m1_n10260_7868# m1_n11408_4493# m1_n11408_4493# m1_n10260_7868#
+ m1_n11408_4493# vdd m1_n11408_4493# vdd m1_n11408_4493# pfet$278
Xpfet$271_7 vdd vdd m1_2446_1478# m1_208_n340# pfet$271
Xnfet$297_7 m1_17703_6956# m1_17703_6956# vss vss m1_18162_6800# vss nfet$297
Xnfet$298_12 m1_15618_7156# vss m1_15755_6960# vss nfet$298
Xnfet$295_4 m1_8596_7868# vss m1_10834_5099# vss nfet$295
Xnfet$293_1 m1_n16410_5099# vss m1_n15874_4493# vss nfet$293
Xpfet$278_1 m1_n6066_7868# m1_n6066_7868# m1_n7214_4493# vdd m1_n7214_4493# m1_n6066_7868#
+ vdd vdd m1_n7214_4493# m1_n6066_7868# m1_n7214_4493# m1_n7214_4493# m1_n6066_7868#
+ m1_n7214_4493# vdd m1_n7214_4493# vdd m1_n7214_4493# pfet$278
Xnfet$298_13 ref vss m1_16242_6960# vss nfet$298
Xnfet$293_2 m1_n12216_5099# vss m1_n11680_4493# vss nfet$293
Xnfet$295_5 m1_4402_7868# vss m1_6640_5099# vss nfet$295
Xpfet$278_2 m1_n14454_7868# m1_n14454_7868# m1_n15602_4493# vdd m1_n15602_4493# m1_n14454_7868#
+ vdd vdd m1_n15602_4493# m1_n14454_7868# m1_n15602_4493# m1_n15602_4493# m1_n14454_7868#
+ m1_n15602_4493# vdd m1_n15602_4493# vdd m1_n15602_4493# pfet$278
Xpfet$283_0 vdd vdd m1_n2336_5099# m1_n4030_5270# pfet$283
Xnfet$295_6 m1_208_n340# vss m1_2446_1478# vss nfet$295
Xpfet$275_10 vdd vdd m1_15618_7156# m1_12790_7868# pfet$275
Xnfet$291_0 m1_3254_n340# vss m1_2982_n340# m1_2982_n340# m1_2982_n340# m1_3254_n340#
+ m1_3254_n340# vss m1_2982_n340# vss nfet$291
Xpfet$276_0 vdd m1_16599_2028# m1_17703_788# m1_15618_394# pfet$276
Xpfet$275_11 vdd vdd m1_16599_5522# m1_15979_5220# pfet$275
Xnfet$295_7 m1_208_7868# vss m1_2446_5099# vss nfet$295
Xpfet$276_1 vdd m1_16242_n208# m1_15979_2344# m1_15755_n208# pfet$276
Xnfet$291_1 m1_7448_n340# vss m1_7176_n340# m1_7176_n340# m1_7176_n340# m1_7448_n340#
+ m1_7448_n340# vss m1_7176_n340# vss nfet$291
Xpfet$275_12 vdd vdd m1_16242_6960# ref pfet$275
Xpfet$276_2 vdd m1_15979_2344# m1_16243_1828# m1_15618_394# pfet$276
Xnfet$291_2 m1_11642_n340# vss m1_11370_n340# m1_11370_n340# m1_11370_n340# m1_11642_n340#
+ m1_11642_n340# vss m1_11370_n340# vss nfet$291
Xpfet$281_0 vdd vdd m1_n8022_5099# m1_n10260_7868# pfet$281
Xpfet$275_13 vdd vdd m1_15755_6960# m1_15618_7156# pfet$275
Xpfet$276_3 vdd m1_17703_788# m1_18496_1828# m1_15755_n208# pfet$276
Xnfet$291_3 m1_n940_n340# vss m1_n1212_n340# m1_n1212_n340# m1_n1212_n340# m1_n940_n340#
+ m1_n940_n340# vss m1_n1212_n340# vss nfet$291
Xpfet$274_0 m1_7448_n340# vdd vdd m1_7448_n340# m1_7176_n340# m1_7176_n340# m1_7448_n340#
+ vdd m1_7176_n340# m1_7176_n340# pfet$274
Xnfet$302_0 m1_19469_4920# m1_19469_4920# m1_19675_2344# m1_19675_2344# m1_19911_1672#
+ vss nfet$302
Xpfet$281_1 vdd vdd m1_n16410_5099# div pfet$281
Xnfet$291_4 m1_11642_4493# vss m1_11370_4493# m1_11370_4493# m1_11370_4493# m1_11642_4493#
+ m1_11642_4493# vss m1_11370_4493# vss nfet$291
Xpfet$276_4 vdd m1_17703_6956# m1_18496_5840# m1_15755_6960# pfet$276
Xpfet$274_1 m1_11642_n340# vdd vdd m1_11642_n340# m1_11370_n340# m1_11370_n340# m1_11642_n340#
+ vdd m1_11370_n340# m1_11370_n340# pfet$274
Xpfet$281_2 vdd vdd m1_n12216_5099# m1_n14454_7868# pfet$281
Xnfet$302_1 m1_19469_1832# m1_19469_1832# vss vss m1_19911_1672# vss nfet$302
Xnfet$291_5 m1_7448_4493# vss m1_7176_4493# m1_7176_4493# m1_7176_4493# m1_7448_4493#
+ m1_7448_4493# vss m1_7176_4493# vss nfet$291
Xpfet$276_5 vdd m1_15979_5220# m1_16243_5840# m1_15618_7156# pfet$276
Xpfet$274_2 m1_3254_n340# vdd vdd m1_3254_n340# m1_2982_n340# m1_2982_n340# m1_3254_n340#
+ vdd m1_2982_n340# m1_2982_n340# pfet$274
Xnfet$291_6 m1_n940_4493# vss m1_n1212_4493# m1_n1212_4493# m1_n1212_4493# m1_n940_4493#
+ m1_n940_4493# vss m1_n1212_4493# vss nfet$291
Xpfet$276_6 vdd m1_16599_5522# m1_17703_6956# m1_15618_7156# pfet$276
Xpfet$272_0 vdd vdd m1_7176_n340# m1_6640_1478# pfet$272
Xpfet$274_3 m1_n940_n340# vdd vdd m1_n940_n340# m1_n1212_n340# m1_n1212_n340# m1_n940_n340#
+ vdd m1_n1212_n340# m1_n1212_n340# pfet$274
.ends

.subckt pfet$311 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=9.75p pd=31.3u as=9.75p ps=31.3u w=15u l=0.5u
.ends

.subckt nfet$330 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.5u
.ends

.subckt pfet$313 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$331 a_n84_0# a_38_n132# a_138_0# VSUBS
X0 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.5u
.ends

.subckt cap_mim$5 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
.ends

.subckt pfet$312 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=9.75p pd=31.3u as=9.75p ps=31.3u w=15u l=0.5u
.ends

.subckt nfet$332 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt CSRVCO_20250823$1 vctrl vosc vdd vss
Xpfet$311_11 vdd m1_n12264_2422# m1_n11916_1270# m1_n9352_266# pfet$311
Xnfet$330_0 m1_n9838_266# m1_n12754_674# m1_n9352_266# vss nfet$330
Xpfet$311_12 vdd m1_n14693_3963# m1_n11296_266# m1_n11782_266# pfet$311
Xnfet$330_1 vctrl vss m1_n12268_985# vss nfet$330
Xpfet$311_13 vdd m1_n13722_3340# m1_n10324_266# m1_n10810_266# pfet$311
Xpfet$311_14 vdd m1_n15180_4275# m1_n11782_266# m1_n11916_1270# pfet$311
Xnfet$330_2 vctrl vss m1_n14283_186# vss nfet$330
Xpfet$313_0 vdd vdd vosc m1_n8380_274# pfet$313
Xnfet$330_3 vctrl vss m1_n13794_186# vss nfet$330
Xpfet$313_1 vdd vdd m1_n8380_274# m1_n11916_1270# pfet$313
Xnfet$330_4 vctrl vss m1_n13240_368# vss nfet$330
Xnfet$330_5 vctrl vss m1_n12754_674# vss nfet$330
Xnfet$330_6 vctrl m1_n16019_266# vss vss nfet$330
Xpfet$311_0 vdd vdd m1_n12264_2422# m1_n16019_266# pfet$311
Xnfet$330_7 vctrl vss m1_n15245_186# vss nfet$330
Xpfet$311_1 vdd vdd m1_n14208_3657# m1_n16019_266# pfet$311
Xnfet$330_8 vctrl vss m1_n14765_186# vss nfet$330
Xpfet$311_2 vdd vdd m1_n13722_3340# m1_n16019_266# pfet$311
Xnfet$330_9 m1_n10324_266# m1_n13240_368# m1_n9838_266# vss nfet$330
Xpfet$311_4 vdd vdd m1_n13236_3035# m1_n16019_266# pfet$311
Xpfet$311_3 vdd m1_n16019_266# vdd m1_n16019_266# pfet$311
Xpfet$311_5 vdd vdd m1_n14693_3963# m1_n16019_266# pfet$311
Xpfet$311_6 vdd vdd m1_n12750_2729# m1_n16019_266# pfet$311
Xpfet$311_7 vdd vdd m1_n15180_4275# m1_n16019_266# pfet$311
Xpfet$311_8 vdd m1_n13236_3035# m1_n9838_266# m1_n10324_266# pfet$311
Xpfet$311_9 vdd m1_n12750_2729# m1_n9352_266# m1_n9838_266# pfet$311
Xnfet$331_0 vss vss vss vss nfet$331
Xnfet$331_1 vss vss vss vss nfet$331
Xnfet$330_10 m1_n9352_266# m1_n12268_985# m1_n11916_1270# vss nfet$330
Xnfet$330_11 m1_n11916_1270# m1_n15245_186# m1_n11782_266# vss nfet$330
Xcap_mim$5_0 vss m1_n11296_266# cap_mim$5
Xnfet$330_12 m1_n11782_266# m1_n14765_186# m1_n11296_266# vss nfet$330
Xcap_mim$5_1 vss m1_n10810_266# cap_mim$5
Xnfet$330_13 m1_n11296_266# m1_n14283_186# m1_n10810_266# vss nfet$330
Xnfet$330_14 m1_n10810_266# m1_n13794_186# m1_n10324_266# vss nfet$330
Xpfet$312_0 vdd vdd vdd vdd pfet$312
Xcap_mim$5_2 vss m1_n10324_266# cap_mim$5
Xcap_mim$5_3 vss m1_n11916_1270# cap_mim$5
Xpfet$312_1 vdd vdd vdd vdd pfet$312
Xcap_mim$5_4 vss m1_n9352_266# cap_mim$5
Xcap_mim$5_5 vss m1_n9838_266# cap_mim$5
Xcap_mim$5_6 vss m1_n11782_266# cap_mim$5
Xnfet$332_0 m1_n8380_274# vss vosc vss nfet$332
Xnfet$332_1 m1_n11916_1270# vss m1_n8380_274# vss nfet$332
Xpfet$311_10 vdd m1_n14208_3657# m1_n10810_266# m1_n11296_266# pfet$311
.ends

.subckt top_level_20250912_nosc i_cp_100u div_def div_prc_s8 div_prc_s7 div_prc_s6
+ div_prc_s5 div_prc_s4 div_prc_s3 div_prc_s2 div_prc_s1 div_prc_s0 div_out div_in
+ div_swc_s0 div_swc_s1 div_swc_s2 div_swc_s3 div_swc_s4 div_swc_s5 div_swc_s6 div_swc_s7
+ div_swc_s8 lock ref ext_pfd_div ext_pfd_ref ext_pfd_up ext_pfd_down mx_pfd_s1 mx_pfd_s0
+ down cp_s1 cp_s2 cp_s3 cp_s4 filter_in filter_out mx_vco_s0 mx_vco_s1 div_rpc_s0
+ div_rsc_s0 div_rsc_s1 div_rpc_s1 div_rsc_s2 div_rpc_s2 div_rsc_s3 div_rsc_s4 div_rsc_s5
+ div_rsc_s6 div_rsc_s7 div_rsc_s8 div_rpc_s3 div_rpc_s4 div_rpc_s5 div_rpc_s6 div_rpc_s7
+ div_rpc_s8 mx_ref_s1 mx_ref_s0 xp_3_1_MUX$2_0/B_1 BIAS$1_0/200n xp_3_1_MUX$2_1/B_1
+ ext_vco_out up vss BIAS$1_0/200p2 BIAS$1_0/200p1 out ext_vco_in vdd
Xasc_hysteresis_buffer$4_0 vss ref vdd xp_3_1_MUX$3_0/OUT_1 asc_hysteresis_buffer$4
Xxp_3_1_MUX$3_1 mx_ref_s0 mx_ref_s1 vdd vss xp_3_1_MUX$3_1/OUT_1 xp_3_1_MUX$3_1/C_1
+ xp_3_1_MUX$3_1/B_1 xp_3_1_MUX$3_1/A_1 xp_3_1_MUX$3
Xxp_3_1_MUX$3_0 mx_ref_s0 mx_ref_s1 vdd vss xp_3_1_MUX$3_0/OUT_1 xp_3_1_MUX$3_1/C_1
+ xp_3_1_MUX$3_0/B_1 xp_3_1_MUX$3_0/A_1 xp_3_1_MUX$3
Xasc_dual_psd_def_20250809$3_0 vdd vss div_rpc_s0 div_rpc_s1 div_rpc_s2 div_rpc_s3
+ div_rpc_s4 div_rpc_s5 div_rpc_s6 div_rpc_s7 div_rpc_s8 xp_3_1_MUX$3_1/B_1 div_rsc_s0
+ div_rsc_s1 div_rsc_s2 div_rsc_s3 div_rsc_s4 div_rsc_s5 div_rsc_s6 div_rsc_s7 div_rsc_s8
+ xp_3_1_MUX$3_0/B_1 vss asc_dual_psd_def_20250809$3
Xasc_drive_buffer$3_0 vss xp_3_1_MUX$2_0/OUT_1 vdd asc_drive_buffer$2_0/in asc_drive_buffer$3
Xasc_hysteresis_buffer$3_0 vss xp_3_1_MUX$3_1/OUT_1 vdd xp_3_1_MUX$2_3/OUT_1 asc_hysteresis_buffer$3
Xxp_3_1_MUX$2_0 mx_vco_s0 mx_vco_s1 vdd vss xp_3_1_MUX$2_0/OUT_1 xp_3_1_MUX$2_0/C_1
+ xp_3_1_MUX$2_0/B_1 ext_vco_out xp_3_1_MUX$2
Xxp_3_1_MUX$2_1 mx_vco_s0 mx_vco_s1 vdd vss filter_out xp_3_1_MUX$2_1/C_1 xp_3_1_MUX$2_1/B_1
+ ext_vco_in xp_3_1_MUX$2
Xxp_3_1_MUX$2_2 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX$2_2/OUT_1 xp_3_1_MUX$2_2/C_1
+ xp_3_1_MUX$2_2/B_1 ext_pfd_up xp_3_1_MUX$2
Xxp_programmable_basic_pump$1_0 asc_drive_buffer_up$1_0/out vdd cp_s1 cp_s2 cp_s3
+ cp_s4 asc_drive_buffer$2_6/out filter_in BIAS$1_0/100n vss xp_programmable_basic_pump$1
Xxp_3_1_MUX$2_4 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX$2_4/OUT_1 xp_3_1_MUX$2_4/C_1
+ xp_3_1_MUX$2_4/B_1 ext_pfd_div xp_3_1_MUX$2
Xxp_3_1_MUX$2_3 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX$2_3/OUT_1 xp_3_1_MUX$2_3/C_1
+ xp_3_1_MUX$2_3/B_1 ext_pfd_ref xp_3_1_MUX$2
Xasc_dual_psd_def_20250809$2_0 vdd vss div_prc_s0 div_prc_s1 div_prc_s2 div_prc_s3
+ div_prc_s4 div_prc_s5 div_prc_s6 div_prc_s7 div_prc_s8 xp_3_1_MUX$2_4/OUT_1 div_swc_s0
+ div_swc_s1 div_swc_s2 div_swc_s3 div_swc_s4 div_swc_s5 div_swc_s6 div_swc_s7 div_swc_s8
+ asc_drive_buffer$2_0/in div_def asc_dual_psd_def_20250809$2
Xxp_3_1_MUX$2_5 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX$2_5/OUT_1 xp_3_1_MUX$2_5/C_1
+ xp_3_1_MUX$2_5/B_1 ext_pfd_down xp_3_1_MUX$2
Xasc_PFD_DFF_20250831$1_0 vss xp_3_1_MUX$2_5/C_1 xp_3_1_MUX$2_2/C_1 vdd xp_3_1_MUX$2_3/C_1
+ xp_3_1_MUX$2_4/C_1 asc_PFD_DFF_20250831$1
Xasc_drive_buffer$2_0 vss asc_drive_buffer$2_0/in vdd div_in asc_drive_buffer$2
Xasc_PFD_DFF_20250831$1_1 vss xp_3_1_MUX$2_2/B_1 xp_3_1_MUX$2_5/B_1 vdd xp_3_1_MUX$2_3/B_1
+ xp_3_1_MUX$2_4/B_1 asc_PFD_DFF_20250831$1
Xasc_drive_buffer$2_1 vss xp_3_1_MUX$2_0/OUT_1 vdd out asc_drive_buffer$2
Xasc_drive_buffer_up$1_0 vss asc_drive_buffer_up$1_0/out xp_3_1_MUX$2_2/OUT_1 vdd
+ asc_drive_buffer_up$1
Xasc_drive_buffer$2_2 vss xp_3_1_MUX$2_4/OUT_1 vdd div_out asc_drive_buffer$2
Xasc_drive_buffer$2_3 vss asc_drive_buffer$2_3/in vdd lock asc_drive_buffer$2
Xasc_drive_buffer$2_4 vss xp_3_1_MUX$2_2/OUT_1 vdd up asc_drive_buffer$2
Xasc_drive_buffer$2_5 vss xp_3_1_MUX$2_5/OUT_1 vdd down asc_drive_buffer$2
Xasc_drive_buffer$2_6 vss xp_3_1_MUX$2_5/OUT_1 vdd asc_drive_buffer$2_6/out asc_drive_buffer$2
XBIAS$1_0 vdd vss BIAS$1_0/100n BIAS$1_0/200n i_cp_100u BIAS$1_0/200p1 BIAS$1_0/200p2
+ BIAS$1
Xasc_lock_detector_20250826$1_0 xp_3_1_MUX$2_3/OUT_1 vdd xp_3_1_MUX$2_4/OUT_1 asc_drive_buffer$2_3/in
+ vss asc_lock_detector_20250826$1
XCSRVCO_20250823$1_0 xp_3_1_MUX$2_1/C_1 xp_3_1_MUX$2_0/C_1 vdd vss CSRVCO_20250823$1
.ends

.subckt nfet$348 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$331 a_750_0# a_546_0# a_446_n60# a_242_n60# w_n180_n88# a_38_n60# a_n92_0#
+ a_342_0# a_138_0# a_650_n60#
X0 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X2 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.5u
.ends

.subckt cap_mim$6 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=50u c_length=100u
.ends

.subckt nfet$346 a_30_n132# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt nfet$351 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.5u
.ends

.subckt ppolyf_u_resistor$4 a_4000_0# a_n376_0# a_n132_0#
X0 a_n132_0# a_4000_0# a_n376_0# ppolyf_u r_width=1u r_length=20u
.ends

.subckt pfet$329 a_28_460# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_460# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt pfet$327 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# w_n180_n88# a_1262_n60# a_38_n60# a_n92_0# a_1058_n60# a_854_n60# a_342_0#
+ a_138_0# a_650_n60# a_1362_0#
X0 a_1362_0# a_1262_n60# a_1158_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X1 a_954_0# a_854_n60# a_750_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X2 a_1566_0# a_1466_n60# a_1362_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.5u
X3 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X4 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X5 a_1158_0# a_1058_n60# a_954_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X6 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.5u
X7 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
.ends

.subckt pfet$332 a_1054_0# a_734_0# a_828_n136# a_28_n136# a_254_0# a_894_0# a_188_n136#
+ a_988_n136# w_n180_n88# a_348_n136# a_1214_0# a_1148_n136# a_414_0# a_n92_0# a_94_0#
+ a_574_0# a_508_n136# a_668_n136#
X0 a_1214_0# a_1148_n136# a_1054_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_734_0# a_668_n136# a_574_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X3 a_574_0# a_508_n136# a_414_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X4 a_1054_0# a_988_n136# a_894_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X5 a_894_0# a_828_n136# a_734_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X6 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X7 a_414_0# a_348_n136# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt pfet$330 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$349 a_750_0# a_546_0# a_446_n132# a_n84_0# a_650_n132# a_38_n132# a_342_0#
+ a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_546_0# a_446_n132# a_342_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X2 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
X3 a_750_0# a_650_n132# a_546_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt nfet$347 a_750_0# a_546_0# a_446_n132# a_n84_0# a_650_n132# a_38_n132# a_342_0#
+ a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.5u
X1 a_546_0# a_446_n132# a_342_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.5u
X2 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.5u
X3 a_750_0# a_650_n132# a_546_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.5u
.ends

.subckt nfet$352 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt nfet$350 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$328 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=0.8125p pd=3.8u as=0.325p ps=1.77u w=1.25u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.325p pd=1.77u as=0.8125p ps=3.8u w=1.25u l=0.5u
.ends

.subckt pfet$325 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_348_n136# a_414_0#
+ a_n92_0# a_94_0# a_574_0# a_508_n136#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_n136# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_n136# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$344 a_254_0# a_30_n132# a_n84_0# a_94_0# a_190_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt nfet$345 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt pfet$326 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
.ends

.subckt OTAforChargePump$2 vdd vss out iref inn inp
Xpfet$325_11 iref vdd iref vdd iref m1_n400_n914# vdd m1_n400_n914# vdd iref pfet$325
Xpfet$325_10 iref vdd iref vdd iref iref vdd iref vdd iref pfet$325
Xnfet$344_0 vss m1_116_n1334# vss out m1_116_n1334# vss nfet$344
Xnfet$344_1 vss m1_116_n1334# vss m1_116_n1334# m1_116_n1334# vss nfet$344
Xnfet$344_2 vss m1_116_n1334# vss m1_116_n1334# m1_116_n1334# vss nfet$344
Xnfet$344_3 vss m1_116_n1334# vss out m1_116_n1334# vss nfet$344
Xpfet$325_0 inn m1_n400_n914# inn vdd inn out m1_n400_n914# out m1_n400_n914# inn
+ pfet$325
Xpfet$325_1 inp m1_n400_n914# inp vdd inp m1_116_n1334# m1_n400_n914# m1_116_n1334#
+ m1_n400_n914# inp pfet$325
Xpfet$325_2 iref vdd iref vdd iref iref vdd iref vdd iref pfet$325
Xpfet$325_3 iref vdd iref vdd iref m1_n400_n914# vdd m1_n400_n914# vdd iref pfet$325
Xpfet$325_5 iref vdd iref vdd iref iref vdd iref vdd iref pfet$325
Xpfet$325_4 iref vdd iref vdd iref m1_n400_n914# vdd m1_n400_n914# vdd iref pfet$325
Xpfet$325_6 iref vdd iref vdd iref iref vdd iref vdd iref pfet$325
Xpfet$325_7 iref vdd iref vdd iref m1_n400_n914# vdd m1_n400_n914# vdd iref pfet$325
Xpfet$325_8 inp m1_n400_n914# inp vdd inp m1_116_n1334# m1_n400_n914# m1_116_n1334#
+ m1_n400_n914# inp pfet$325
Xpfet$325_9 inn m1_n400_n914# inn vdd inn out m1_n400_n914# out m1_n400_n914# inn
+ pfet$325
Xnfet$345_0 vss vss vss vss vss vss vss vss vss vss nfet$345
Xnfet$345_1 vss vss vss vss vss vss vss vss vss vss nfet$345
Xpfet$326_0 m1_n400_n914# m1_n400_n914# m1_n400_n914# vdd m1_n400_n914# m1_n400_n914#
+ pfet$326
Xpfet$326_2 vdd vdd vdd vdd vdd vdd pfet$326
Xpfet$326_1 m1_n400_n914# m1_n400_n914# m1_n400_n914# vdd m1_n400_n914# m1_n400_n914#
+ pfet$326
Xpfet$326_3 vdd vdd vdd vdd vdd vdd pfet$326
Xpfet$326_4 vdd vdd vdd vdd vdd vdd pfet$326
Xpfet$326_5 vdd vdd vdd vdd vdd vdd pfet$326
.ends

.subckt PCP1248X$1 vdd s3 s2 s1 s0 vin iref200u out up down vss
Xnfet$348_0 vss vss vss vss vss vss nfet$348
Xpfet$331_5 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$331
Xcap_mim$6_0 m1_n1751_n2187# vdd cap_mim$6
Xnfet$348_1 vss vss vss vss vss vss nfet$348
Xpfet$331_6 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$331
Xcap_mim$6_1 vss m1_9963_14448# cap_mim$6
Xnfet$348_2 vss m1_9963_14448# vss m1_9963_14448# m1_9963_14448# vss nfet$348
Xpfet$331_7 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$331
Xcap_mim$6_2 vss OTAforChargePump$2_0/out cap_mim$6
Xpfet$331_8 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$331
Xnfet$346_0 s0 m1_n47_11059# m1_1641_5849# vss nfet$346
Xnfet$346_1 s1 m1_n47_11059# m1_n91_6229# vss nfet$346
Xpfet$331_9 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$331
Xnfet$346_2 s3 m1_n47_11059# m1_n1771_4009# vss nfet$346
Xnfet$351_0 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$351
Xnfet$346_3 s2 m1_n47_11059# m1_1137_12199# vss nfet$346
Xppolyf_u_resistor$4_0 m1_3630_13790# vss m1_n502_13390# ppolyf_u_resistor$4
Xpfet$329_0 s0 vdd m1_1641_5849# vdd pfet$329
Xnfet$351_1 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$351
Xnfet$346_4 m1_n539_12403# m1_16753_5552# vss vss nfet$346
Xppolyf_u_resistor$4_1 OTAforChargePump$2_0/inp vss m1_n502_13390# ppolyf_u_resistor$4
Xnfet$351_2 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$351
Xpfet$329_1 s3 vdd m1_n1771_4009# vdd pfet$329
Xnfet$346_5 s0 OTAforChargePump$2_0/out m1_16753_5552# vss nfet$346
Xppolyf_u_resistor$4_2 m1_3630_14590# vss m1_n502_14190# ppolyf_u_resistor$4
Xnfet$351_10 vss vss vss vss vss vss nfet$351
Xpfet$329_2 m1_n1311_12403# vdd m1_n47_11059# m1_n91_6229# pfet$329
Xnfet$351_3 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$351
Xnfet$346_10 m1_n2855_12403# m1_14137_3830# vss vss nfet$346
Xnfet$346_6 m1_n1311_12403# m1_15009_5932# vss vss nfet$346
Xppolyf_u_resistor$4_3 m1_3630_13790# vss m1_n502_14190# ppolyf_u_resistor$4
Xnfet$346_11 s3 OTAforChargePump$2_0/out m1_14137_3830# vss nfet$346
Xnfet$351_11 vss vss vss vss vss vss nfet$351
Xpfet$329_3 m1_n2083_12403# vdd m1_n47_11059# m1_1137_12199# pfet$329
Xpfet$327_0 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$327
Xnfet$351_4 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$351
Xnfet$346_7 s1 OTAforChargePump$2_0/out m1_15009_5932# vss nfet$346
Xppolyf_u_resistor$4_4 m1_3630_14590# vss m1_n502_14990# ppolyf_u_resistor$4
Xpfet$329_4 m1_n2855_12403# vdd m1_n47_11059# m1_n1771_4009# pfet$329
Xnfet$351_5 m1_n47_11059# m1_n47_11059# m1_n47_11059# m1_n47_11059# m1_n47_11059#
+ vss nfet$351
Xpfet$327_1 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$327
Xnfet$346_8 m1_n2083_12403# m1_15881_3450# vss vss nfet$346
Xppolyf_u_resistor$4_5 vdd vss m1_n502_14990# ppolyf_u_resistor$4
Xnfet$351_6 vss vss vss vss vss vss nfet$351
Xpfet$329_5 s1 vdd m1_n91_6229# vdd pfet$329
Xpfet$327_2 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$327
Xpfet$332_0 m1_n2925_n36# m1_n2925_n36# up up out out up up vdd up out up m1_n2925_n36#
+ out m1_n2925_n36# out up up pfet$332
Xnfet$346_9 s2 OTAforChargePump$2_0/out m1_15881_3450# vss nfet$346
Xnfet$351_7 vss vss vss vss vss vss nfet$351
Xpfet$329_6 s2 vdd m1_1137_12199# vdd pfet$329
Xpfet$327_3 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$327
Xpfet$331_10 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$331
Xnfet$351_8 vss vss vss vss vss vss nfet$351
Xpfet$329_7 m1_n539_12403# vdd m1_n47_11059# m1_1641_5849# pfet$329
Xpfet$329_10 m1_n2083_12403# vdd OTAforChargePump$2_0/out m1_15881_3450# pfet$329
Xpfet$327_4 m1_n2925_n36# m1_n2925_n36# m1_n25_493# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n25_493# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36#
+ m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n25_493# m1_n1751_n2187# m1_n25_493#
+ pfet$327
Xpfet$331_11 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$331
Xpfet$329_8 m1_n539_12403# vdd OTAforChargePump$2_0/out m1_16753_5552# pfet$329
Xnfet$351_9 vss vss vss vss vss vss nfet$351
Xpfet$327_5 m1_n47_11059# m1_n47_11059# m1_6759_7857# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n47_11059# m1_6759_7857# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n47_11059# m1_n1751_n2187# m1_n1751_n2187# m1_n47_11059# m1_6759_7857# m1_n1751_n2187#
+ m1_6759_7857# pfet$327
Xpfet$329_11 m1_n2855_12403# vdd OTAforChargePump$2_0/out m1_14137_3830# pfet$329
Xpfet$330_0 vdd vdd m1_n2855_12403# s3 pfet$330
Xpfet$329_9 m1_n1311_12403# vdd OTAforChargePump$2_0/out m1_15009_5932# pfet$329
Xpfet$327_6 vdd vdd m1_6759_7857# m1_n47_11059# m1_n47_11059# vdd m1_6759_7857# m1_n47_11059#
+ vdd m1_n47_11059# m1_n47_11059# vdd m1_n47_11059# m1_n47_11059# vdd m1_6759_7857#
+ m1_n47_11059# m1_6759_7857# pfet$327
Xpfet$330_1 vdd vdd m1_n2083_12403# s2 pfet$330
Xnfet$349_0 vss m1_9475_12045# OTAforChargePump$2_0/out vss OTAforChargePump$2_0/out
+ OTAforChargePump$2_0/out vss m1_9475_12045# OTAforChargePump$2_0/out vss nfet$349
Xpfet$327_7 vdd vdd m1_n25_493# m1_n91_6229# m1_n91_6229# vdd m1_n25_493# m1_n91_6229#
+ vdd m1_n91_6229# m1_n91_6229# vdd m1_n91_6229# m1_n91_6229# vdd m1_n25_493# m1_n91_6229#
+ m1_n25_493# pfet$327
Xpfet$330_2 vdd vdd m1_n539_12403# s0 pfet$330
Xnfet$349_1 vss m1_n1751_n2187# OTAforChargePump$2_0/out vss OTAforChargePump$2_0/out
+ OTAforChargePump$2_0/out vss m1_n1751_n2187# OTAforChargePump$2_0/out vss nfet$349
Xpfet$327_8 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$327
Xpfet$330_3 vdd vdd m1_n1311_12403# s1 pfet$330
Xnfet$349_2 vss m1_9475_12045# OTAforChargePump$2_0/out vss OTAforChargePump$2_0/out
+ OTAforChargePump$2_0/out vss m1_9475_12045# OTAforChargePump$2_0/out vss nfet$349
Xpfet$327_9 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$327
Xnfet$347_30 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$347
Xnfet$349_3 vss m1_n1751_n2187# OTAforChargePump$2_0/out vss OTAforChargePump$2_0/out
+ OTAforChargePump$2_0/out vss m1_n1751_n2187# OTAforChargePump$2_0/out vss nfet$349
Xnfet$347_0 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$347
Xnfet$347_20 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$347
Xnfet$347_31 m1_n47_11059# m1_14015_1164# m1_9963_14448# m1_n47_11059# m1_9963_14448#
+ m1_9963_14448# m1_n47_11059# m1_14015_1164# m1_9963_14448# vss nfet$347
Xnfet$347_1 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$347
Xnfet$347_21 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$347
Xnfet$347_32 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$347
Xnfet$347_10 m1_13543_n1758# m1_15911_n1318# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15911_n1318# m1_9963_14448# vss nfet$347
Xnfet$347_2 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$347
Xnfet$347_22 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$347
Xnfet$347_33 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$347
Xnfet$352_0 down out m1_13543_n1758# down out m1_13543_n1758# down out down vss nfet$352
Xnfet$347_11 m1_13543_n1758# m1_15039_784# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15039_784# m1_9963_14448# vss nfet$347
Xnfet$347_34 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$347
Xnfet$347_23 vss m1_15039_784# m1_15009_5932# vss m1_15009_5932# m1_15009_5932# vss
+ m1_15039_784# m1_15009_5932# vss nfet$347
Xnfet$347_3 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# vss nfet$347
Xnfet$347_12 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$347
Xpfet$327_30 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ pfet$327
Xnfet$347_4 m1_13543_n1758# m1_15039_784# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15039_784# m1_9963_14448# vss nfet$347
Xnfet$347_24 vss vss vss vss vss vss vss vss vss vss nfet$347
Xnfet$347_35 vss m1_14015_1164# OTAforChargePump$2_0/out vss OTAforChargePump$2_0/out
+ OTAforChargePump$2_0/out vss m1_14015_1164# OTAforChargePump$2_0/out vss nfet$347
Xnfet$347_13 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$347
Xpfet$327_31 m1_n2925_n36# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187#
+ m1_1671_n1319# pfet$327
Xpfet$327_20 m1_n2925_n36# m1_n2925_n36# m1_1671_873# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_873# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36#
+ m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_873# m1_n1751_n2187# m1_1671_873#
+ pfet$327
Xnfet$347_36 OTAforChargePump$2_0/inp m1_9475_12045# m1_9963_14448# OTAforChargePump$2_0/inp
+ m1_9963_14448# m1_9963_14448# OTAforChargePump$2_0/inp m1_9475_12045# m1_9963_14448#
+ vss nfet$347
Xnfet$347_25 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$347
Xnfet$347_5 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# vss nfet$347
Xnfet$347_14 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$347
Xnfet$350_0 s3 vss m1_n2855_12403# vss nfet$350
Xpfet$327_10 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$327
Xpfet$327_32 m1_n2925_n36# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187#
+ m1_1671_n1319# pfet$327
Xpfet$327_21 vdd vdd m1_1671_873# m1_1641_5849# m1_1641_5849# vdd m1_1671_873# m1_1641_5849#
+ vdd m1_1641_5849# m1_1641_5849# vdd m1_1641_5849# m1_1641_5849# vdd m1_1671_873#
+ m1_1641_5849# m1_1671_873# pfet$327
Xnfet$347_6 m1_13543_n1758# m1_16783_404# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_16783_404# m1_9963_14448# vss nfet$347
Xnfet$347_26 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$347
Xnfet$347_15 vss vss vss vss vss vss vss vss vss vss nfet$347
Xpfet$328_0 vdd vdd vdd vdd vdd vdd pfet$328
Xnfet$350_1 s2 vss m1_n2083_12403# vss nfet$350
Xpfet$327_11 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$327
Xpfet$327_22 vdd vdd m1_1671_n1319# m1_1137_12199# m1_1137_12199# vdd m1_1671_n1319#
+ m1_1137_12199# vdd m1_1137_12199# m1_1137_12199# vdd m1_1137_12199# m1_1137_12199#
+ vdd m1_1671_n1319# m1_1137_12199# m1_1671_n1319# pfet$327
Xpfet$327_33 vdd vdd m1_1671_n1319# m1_1137_12199# m1_1137_12199# vdd m1_1671_n1319#
+ m1_1137_12199# vdd m1_1137_12199# m1_1137_12199# vdd m1_1137_12199# m1_1137_12199#
+ vdd m1_1671_n1319# m1_1137_12199# m1_1671_n1319# pfet$327
Xnfet$347_27 vss m1_15911_n1318# m1_15881_3450# vss m1_15881_3450# m1_15881_3450#
+ vss m1_15911_n1318# m1_15881_3450# vss nfet$347
Xnfet$347_16 vss m1_16783_404# m1_16753_5552# vss m1_16753_5552# m1_16753_5552# vss
+ m1_16783_404# m1_16753_5552# vss nfet$347
Xnfet$347_7 m1_13543_n1758# m1_15911_n1318# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15911_n1318# m1_9963_14448# vss nfet$347
Xpfet$328_1 vdd vdd vdd m1_n1751_n2187# m1_n1751_n2187# m1_n1751_n2187# pfet$328
Xnfet$350_2 s1 vss m1_n1311_12403# vss nfet$350
Xpfet$327_12 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$327
Xpfet$327_23 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$327
Xpfet$327_34 vdd vdd m1_1671_n1319# m1_1137_12199# m1_1137_12199# vdd m1_1671_n1319#
+ m1_1137_12199# vdd m1_1137_12199# m1_1137_12199# vdd m1_1137_12199# m1_1137_12199#
+ vdd m1_1671_n1319# m1_1137_12199# m1_1671_n1319# pfet$327
Xnfet$347_8 m1_13543_n1758# m1_15911_n1318# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15911_n1318# m1_9963_14448# vss nfet$347
Xnfet$347_28 vss m1_15911_n1318# m1_15881_3450# vss m1_15881_3450# m1_15881_3450#
+ vss m1_15911_n1318# m1_15881_3450# vss nfet$347
Xnfet$347_17 vss m1_15039_784# m1_15009_5932# vss m1_15009_5932# m1_15009_5932# vss
+ m1_15039_784# m1_15009_5932# vss nfet$347
Xpfet$328_2 vdd vdd vdd m1_9963_14448# m1_n1751_n2187# m1_n1751_n2187# pfet$328
Xnfet$350_3 s0 vss m1_n539_12403# vss nfet$350
Xpfet$327_13 m1_n2925_n36# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187#
+ m1_1671_n1319# pfet$327
Xpfet$327_24 vdd vdd m1_n25_493# m1_n91_6229# m1_n91_6229# vdd m1_n25_493# m1_n91_6229#
+ vdd m1_n91_6229# m1_n91_6229# vdd m1_n91_6229# m1_n91_6229# vdd m1_n25_493# m1_n91_6229#
+ m1_n25_493# pfet$327
Xpfet$327_35 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ pfet$327
XOTAforChargePump$2_0 vdd vss OTAforChargePump$2_0/out iref200u vin OTAforChargePump$2_0/inp
+ OTAforChargePump$2
Xnfet$347_9 m1_13543_n1758# m1_15911_n1318# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15911_n1318# m1_9963_14448# vss nfet$347
Xpfet$328_3 vdd vdd vdd m1_n1751_n2187# m1_n1751_n2187# m1_n1751_n2187# pfet$328
Xnfet$347_29 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$347
Xnfet$347_18 vss m1_15911_n1318# m1_15881_3450# vss m1_15881_3450# m1_15881_3450#
+ vss m1_15911_n1318# m1_15881_3450# vss nfet$347
Xpfet$327_14 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$327
Xpfet$327_25 vdd vdd m1_1671_n1319# m1_1137_12199# m1_1137_12199# vdd m1_1671_n1319#
+ m1_1137_12199# vdd m1_1137_12199# m1_1137_12199# vdd m1_1137_12199# m1_1137_12199#
+ vdd m1_1671_n1319# m1_1137_12199# m1_1671_n1319# pfet$327
Xnfet$347_19 vss m1_15911_n1318# m1_15881_3450# vss m1_15881_3450# m1_15881_3450#
+ vss m1_15911_n1318# m1_15881_3450# vss nfet$347
Xpfet$328_4 vdd vdd vdd m1_9963_14448# m1_n1751_n2187# m1_n1751_n2187# pfet$328
Xpfet$327_15 m1_n2925_n36# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187#
+ m1_1671_n1319# pfet$327
Xpfet$327_26 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$327
Xpfet$328_5 vdd vdd vdd vdd vdd vdd pfet$328
Xpfet$327_16 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ pfet$327
Xpfet$327_27 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$327
Xpfet$331_0 m1_n47_11059# m1_n47_11059# m1_n47_11059# m1_n47_11059# vdd m1_n47_11059#
+ m1_n47_11059# m1_n47_11059# m1_n47_11059# m1_n47_11059# pfet$331
Xpfet$327_17 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$327
Xpfet$327_28 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$327
Xpfet$331_1 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$331
Xpfet$327_18 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$327
Xpfet$327_29 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ pfet$327
Xpfet$331_2 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$331
Xpfet$331_3 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$331
Xpfet$327_19 m1_n2925_n36# m1_n2925_n36# m1_n25_493# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n25_493# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36#
+ m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n25_493# m1_n1751_n2187# m1_n25_493#
+ pfet$327
Xpfet$331_4 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$331
.ends

.subckt pfet$341 a_28_460# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_460# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt nfet$361 a_n84_0# a_94_0# a_30_460# VSUBS
X0 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$340 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=2.6p pd=9.3u as=2.6p ps=9.3u w=4u l=0.28u
.ends

.subckt nfet$362 a_30_n132# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt SCHMITT$3 VDD VSS IN OUT
Xpfet$341_0 OUT VDD m1_596_1544# VSS pfet$341
Xnfet$361_0 m1_592_402# OUT IN VSS nfet$361
Xnfet$361_1 VSS m1_592_402# IN VSS nfet$361
Xpfet$340_0 IN VDD m1_596_1544# OUT pfet$340
Xpfet$340_1 IN VDD VDD m1_596_1544# pfet$340
Xnfet$362_0 OUT m1_592_402# VDD VSS nfet$362
.ends

.subckt nfet$353 a_n84_0# a_94_0# a_30_160# VSUBS
X0 a_94_0# a_30_160# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.28u
.ends

.subckt pfet$333 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt SRLATCH vdd vss q qb s r
Xnfet$353_0 vss qb r vss nfet$353
Xnfet$353_2 q vss s vss nfet$353
Xnfet$353_1 vss qb q vss nfet$353
Xnfet$353_3 q vss qb vss nfet$353
Xpfet$333_0 r vdd m1_818_875# qb pfet$333
Xpfet$333_1 q vdd vdd m1_818_875# pfet$333
Xpfet$333_3 qb vdd q m1_50_875# pfet$333
Xpfet$333_2 s vdd m1_50_875# vdd pfet$333
.ends

.subckt nfet$363 a_30_260# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_260# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt cap_mim$7 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=60u c_length=100u
.ends

.subckt ppolyf_u_resistor$5 a_n376_0# a_4200_0# a_n132_0#
X0 a_n132_0# a_4200_0# a_n376_0# ppolyf_u r_width=1u r_length=21u
.ends

.subckt pfet$342 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt pfet$336 a_254_0# a_348_560# w_n180_n88# a_414_0# a_n92_0# a_94_0# a_574_0#
+ a_508_560# a_188_560# a_28_560#
X0 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt pfet$334 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_348_n136# a_414_0#
+ a_n92_0# a_94_0# a_574_0# a_508_n136#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_n136# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_n136# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$356 a_254_0# a_350_460# a_414_0# a_n84_0# a_94_0# a_510_460# a_190_460#
+ a_574_0# a_30_460# VSUBS
X0 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_460# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_460# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt nfet$354 a_254_0# a_n84_0# a_94_0# a_190_460# a_30_460# VSUBS
X0 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$335 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
.ends

.subckt nfet$357 a_n84_0# a_94_0# a_30_460# VSUBS
X0 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt nfet$355 a_1054_0# a_734_0# a_254_0# a_350_460# a_830_460# a_894_0# a_990_460#
+ a_1214_0# a_414_0# a_n84_0# a_94_0# a_510_460# a_190_460# a_574_0# a_670_460# a_1150_460#
+ a_30_460# VSUBS
X0 a_734_0# a_670_460# a_574_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_574_0# a_510_460# a_414_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X3 a_1054_0# a_990_460# a_894_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X4 a_894_0# a_830_460# a_734_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X5 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X6 a_414_0# a_350_460# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X7 a_1214_0# a_1150_460# a_1054_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt Ncomparator$1 iref vss vdd out inn inp
Xpfet$336_1 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$336
Xpfet$336_0 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$336
Xpfet$336_2 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$336
Xpfet$334_0 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_570_1653# vdd m1_570_1653#
+ vdd m1_1242_549# pfet$334
Xpfet$336_3 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$336
Xpfet$334_1 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_1242_549# vdd m1_1242_549#
+ vdd m1_1242_549# pfet$334
Xpfet$334_2 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_570_1653# vdd m1_570_1653#
+ vdd m1_1242_549# pfet$334
Xpfet$334_3 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_1242_549# vdd m1_1242_549#
+ vdd m1_1242_549# pfet$334
Xnfet$356_0 vss iref m1_506_n191# vss m1_506_n191# iref iref vss iref vss nfet$356
Xnfet$356_1 vss iref iref vss iref iref iref vss iref vss nfet$356
Xnfet$356_2 m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191#
+ m1_506_n191# m1_506_n191# m1_506_n191# vss nfet$356
Xnfet$356_3 m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191#
+ m1_506_n191# m1_506_n191# m1_506_n191# vss nfet$356
Xnfet$354_0 m1_506_n191# m1_506_n191# m1_570_1653# inp inp vss nfet$354
Xnfet$356_4 vss iref iref vss iref iref iref vss iref vss nfet$356
Xnfet$354_1 m1_506_n191# m1_506_n191# m1_1242_549# inn inn vss nfet$354
Xnfet$354_2 m1_506_n191# m1_506_n191# m1_570_1653# inp inp vss nfet$354
Xnfet$356_5 vss iref m1_506_n191# vss m1_506_n191# iref iref vss iref vss nfet$356
Xnfet$354_3 m1_506_n191# m1_506_n191# m1_1242_549# inn inn vss nfet$354
Xpfet$335_0 vdd vdd vdd vdd vdd vdd pfet$335
Xpfet$335_1 vdd vdd vdd vdd vdd vdd pfet$335
Xpfet$335_2 vdd vdd vdd vdd vdd vdd pfet$335
Xpfet$335_3 vdd vdd vdd vdd vdd vdd pfet$335
Xnfet$357_0 vss vss vss vss nfet$357
Xnfet$357_1 vss vss vss vss nfet$357
Xnfet$355_0 out out vss iref iref vss iref vss out vss out iref iref vss iref iref
+ iref vss nfet$355
.ends

.subckt nfet$360 a_254_0# a_n84_0# a_94_0# a_190_460# a_30_460# VSUBS
X0 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$338 a_254_0# a_348_560# w_n180_n88# a_414_0# a_n92_0# a_94_0# a_574_0#
+ a_508_560# a_188_560# a_28_560#
X0 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$358 a_1054_0# a_734_0# a_510_n132# a_254_0# a_894_0# a_670_n132# a_1214_0#
+ a_830_n132# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132# a_574_0# a_990_n132#
+ a_350_n132# a_1150_n132# VSUBS
X0 a_734_0# a_670_n132# a_574_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X3 a_1054_0# a_990_n132# a_894_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X4 a_894_0# a_830_n132# a_734_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X5 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X6 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X7 a_1214_0# a_1150_n132# a_1054_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt pfet$339 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=1.625p ps=6.3u w=2.5u l=0.28u
.ends

.subckt pfet$337 a_1054_0# a_734_0# a_254_0# a_894_0# a_348_560# a_828_560# a_988_560#
+ w_n180_n88# a_1214_0# a_414_0# a_n92_0# a_94_0# a_574_0# a_508_560# a_188_560# a_668_560#
+ a_1148_560# a_28_560#
X0 a_1214_0# a_1148_560# a_1054_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_734_0# a_668_560# a_574_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X3 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X4 a_1054_0# a_988_560# a_894_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X5 a_894_0# a_828_560# a_734_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X6 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X7 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$359 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt Pcomparator$1 vss vdd out iref inn inp
Xnfet$360_0 vss vss m1_3615_n1223# m1_3615_n1223# m1_3615_n1223# vss nfet$360
Xnfet$360_1 vss vss m1_5539_n2811# m1_3615_n1223# m1_3615_n1223# vss nfet$360
Xpfet$338_0 m1_2779_n1752# inp vdd m1_5539_n2811# m1_2779_n1752# m1_5539_n2811# m1_2779_n1752#
+ inp inp inp pfet$338
Xpfet$338_2 m1_2779_n1752# inn vdd m1_3615_n1223# m1_2779_n1752# m1_3615_n1223# m1_2779_n1752#
+ inn inn inn pfet$338
Xnfet$360_3 vss vss m1_3615_n1223# m1_3615_n1223# m1_3615_n1223# vss nfet$360
Xnfet$360_2 vss vss m1_5539_n2811# m1_3615_n1223# m1_3615_n1223# vss nfet$360
Xpfet$338_1 m1_2779_n1752# m1_2779_n1752# vdd m1_2779_n1752# m1_2779_n1752# m1_2779_n1752#
+ m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# pfet$338
Xpfet$338_3 m1_2779_n1752# m1_2779_n1752# vdd m1_2779_n1752# m1_2779_n1752# m1_2779_n1752#
+ m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# pfet$338
Xpfet$338_4 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$338
Xpfet$338_5 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$338
Xpfet$338_6 vdd iref vdd iref vdd iref vdd iref iref iref pfet$338
Xpfet$338_7 vdd iref vdd iref vdd iref vdd iref iref iref pfet$338
Xpfet$338_8 vdd iref vdd iref vdd iref vdd iref iref iref pfet$338
Xpfet$338_9 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$338
Xnfet$358_0 out out m1_5539_n2811# vss vss m1_5539_n2811# vss m1_5539_n2811# out m1_5539_n2811#
+ vss out m1_5539_n2811# vss m1_5539_n2811# m1_5539_n2811# m1_5539_n2811# vss nfet$358
Xpfet$339_0 vdd vdd vdd vdd pfet$339
Xpfet$339_1 vdd vdd vdd vdd pfet$339
Xpfet$339_2 vdd vdd vdd vdd pfet$339
Xpfet$337_0 out out vdd vdd iref iref iref vdd vdd out vdd out vdd iref iref iref
+ iref iref pfet$337
Xpfet$339_3 vdd vdd vdd vdd pfet$339
Xpfet$337_1 out out vdd vdd iref iref iref vdd vdd out vdd out vdd iref iref iref
+ iref iref pfet$337
Xpfet$338_10 vdd iref vdd iref vdd iref vdd iref iref iref pfet$338
Xpfet$338_11 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$338
Xpfet$338_12 m1_2779_n1752# inn vdd m1_3615_n1223# m1_2779_n1752# m1_3615_n1223# m1_2779_n1752#
+ inn inn inn pfet$338
Xnfet$359_0 vss vss vss vss vss vss vss vss vss vss nfet$359
Xpfet$338_13 m1_2779_n1752# inp vdd m1_5539_n2811# m1_2779_n1752# m1_5539_n2811# m1_2779_n1752#
+ inp inp inp pfet$338
Xnfet$359_1 vss vss vss vss vss vss vss vss vss vss nfet$359
.ends

.subckt VCOfinal s3 s0 s1 s2 iref200 fout foutb vss irefn irefp vin a_11641_n18839#
+ vdd
XPCP1248X$1_0 vdd s3 s2 s1 s0 vin iref200 PCP1248X$1_0/out PCP1248X$1_0/up SRLATCH_0/qb
+ vss PCP1248X$1
XSCHMITT$3_1 vdd vss SRLATCH_0/q SCHMITT$3_1/OUT SCHMITT$3
XSRLATCH_0 vdd vss SRLATCH_0/q SRLATCH_0/qb SRLATCH_0/s SRLATCH_0/r SRLATCH
Xnfet$363_0 SRLATCH_0/q vss PCP1248X$1_0/up vss nfet$363
Xnfet$363_1 SCHMITT$3_0/OUT vss foutb vss nfet$363
Xnfet$363_2 SCHMITT$3_1/OUT vss fout vss nfet$363
Xcap_mim$7_0 vss PCP1248X$1_0/out cap_mim$7
Xppolyf_u_resistor$5_0 vss vss Pcomparator$1_0/inp ppolyf_u_resistor$5
Xpfet$342_0 SRLATCH_0/q vdd vdd PCP1248X$1_0/up pfet$342
Xppolyf_u_resistor$5_1 vss m1_13996_n13334# Ncomparator$1_0/inn ppolyf_u_resistor$5
Xpfet$342_1 SCHMITT$3_0/OUT vdd vdd foutb pfet$342
Xppolyf_u_resistor$5_2 vss m1_13996_n13334# Pcomparator$1_0/inp ppolyf_u_resistor$5
Xppolyf_u_resistor$5_3 vss vdd Ncomparator$1_0/inn ppolyf_u_resistor$5
Xpfet$342_2 SCHMITT$3_1/OUT vdd vdd fout pfet$342
XNcomparator$1_0 irefn vss vdd SRLATCH_0/s Ncomparator$1_0/inn PCP1248X$1_0/out Ncomparator$1
XSCHMITT$3_0 vdd vss SRLATCH_0/qb SCHMITT$3_0/OUT SCHMITT$3
XPcomparator$1_0 vss vdd SRLATCH_0/r irefp PCP1248X$1_0/out Pcomparator$1_0/inp Pcomparator$1
.ends

.subckt pfet$322 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt nfet$342 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$340 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt pfet$323 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$321 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt nfet$343 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$341 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt pfet$324 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt qw_NOLclk$1 CLK VDDd VSSd PHI_1 PHI_2
Xpfet$322_1 m1_15103_233# VDDd VDDd m1_13930_233# pfet$322
Xpfet$322_2 m1_12351_431# VDDd VDDd m1_15103_1818# pfet$322
Xpfet$322_3 m1_15103_1818# VDDd VDDd m1_13930_1818# pfet$322
Xnfet$342_0 m1_11601_71# VSSd PHI_1 VSSd nfet$342
Xnfet$342_1 m1_11161_409# VSSd m1_11379_n171# VSSd nfet$342
Xnfet$342_2 m1_11601_2380# VSSd PHI_2 VSSd nfet$342
Xnfet$342_3 CLK VSSd m1_11161_409# VSSd nfet$342
Xnfet$340_0 PHI_1 VSSd m1_13930_233# VSSd nfet$340
Xnfet$340_1 PHI_2 VSSd m1_13930_1818# VSSd nfet$340
Xpfet$323_0 VDDd VDDd PHI_1 m1_11601_71# pfet$323
Xpfet$323_1 VDDd VDDd m1_11379_n171# m1_11161_409# pfet$323
Xpfet$323_2 VDDd VDDd PHI_2 m1_11601_2380# pfet$323
Xpfet$323_3 VDDd VDDd m1_11161_409# CLK pfet$323
Xpfet$321_0 VDDd VDDd m1_13930_233# PHI_1 pfet$321
Xpfet$321_1 VDDd VDDd m1_13930_1818# PHI_2 pfet$321
Xnfet$343_0 m1_12351_431# m1_12351_431# m1_11601_71# m1_11601_71# m1_11837_749# VSSd
+ nfet$343
Xnfet$343_1 m1_11379_n171# m1_11379_n171# VSSd VSSd m1_11837_749# VSSd nfet$343
Xnfet$343_2 m1_12351_2064# m1_12351_2064# m1_11601_2380# m1_11601_2380# m1_11837_1708#
+ VSSd nfet$343
Xnfet$343_3 m1_11161_409# m1_11161_409# VSSd VSSd m1_11837_1708# VSSd nfet$343
Xnfet$341_0 m1_12351_2064# m1_15103_233# VSSd VSSd nfet$341
Xnfet$341_1 m1_15103_233# m1_13930_233# VSSd VSSd nfet$341
Xnfet$341_2 m1_12351_431# m1_15103_1818# VSSd VSSd nfet$341
Xnfet$341_3 m1_15103_1818# m1_13930_1818# VSSd VSSd nfet$341
Xpfet$324_0 VDDd m1_11601_71# VDDd m1_11379_n171# pfet$324
Xpfet$324_1 VDDd VDDd m1_11601_71# m1_12351_431# pfet$324
Xpfet$324_2 VDDd m1_11601_2380# VDDd m1_11161_409# pfet$324
Xpfet$324_3 VDDd VDDd m1_11601_2380# m1_12351_2064# pfet$324
Xpfet$322_0 m1_12351_2064# VDDd VDDd m1_15103_233# pfet$322
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__latq_1$4 D E Q VDD VSS VNW VPW
X0 VSS a_1020_652# Q VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X1 a_504_110# a_36_92# VDD VNW pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X2 VDD a_1020_652# Q VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X3 a_1264_107# a_36_92# a_1020_652# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X4 VSS E a_36_92# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X5 VSS a_1364_532# a_1264_107# VPW nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X6 VDD E a_36_92# VNW pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X7 VDD a_1364_532# a_1224_652# VNW pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X8 a_872_652# D VDD VNW pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X9 a_1364_532# a_1020_652# VDD VNW pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X10 a_1020_652# a_504_110# a_872_107# VPW nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X11 a_872_107# D VSS VPW nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X12 a_1020_652# a_36_92# a_872_652# VNW pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X13 a_504_110# a_36_92# VSS VPW nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X14 a_1364_532# a_1020_652# VSS VPW nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X15 a_1224_652# a_504_110# a_1020_652# VNW pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt DFF_2phase_1$3 VDDd D Q PHI_1 PHI_2 VSSd
Xgf180mcu_fd_sc_mcu9t5v0__latq_1$4_1 D PHI_1 gf180mcu_fd_sc_mcu9t5v0__latq_1$4_1/Q
+ VDDd VSSd VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1$4
Xgf180mcu_fd_sc_mcu9t5v0__latq_1$4_0 gf180mcu_fd_sc_mcu9t5v0__latq_1$4_1/Q PHI_2 Q
+ VDDd VSSd VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1$4
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1$3 I VDD VSS ZN VNW VPW
X0 ZN I VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__and2_1$3 A1 A2 VDD VSS Z VNW VPW
X0 VDD A2 a_36_201# VNW pfet_05v0 ad=0.5054p pd=2.57u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1 a_244_201# A1 a_36_201# VPW nfet_05v0 ad=0.1056p pd=0.98u as=0.2904p ps=2.2u w=0.66u l=0.6u
X2 Z a_36_201# VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.3894p ps=2.06u w=1.32u l=0.6u
X3 Z a_36_201# VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.5054p ps=2.57u w=1.83u l=0.5u
X4 VSS A2 a_244_201# VPW nfet_05v0 ad=0.3894p pd=2.06u as=0.1056p ps=0.98u w=0.66u l=0.6u
X5 a_36_201# A1 VDD VNW pfet_05v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__or2_1$3 A1 A2 VDD VSS Z VNW VPW
X0 a_255_756# A1 a_67_756# VNW pfet_05v0 ad=0.2379p pd=1.435u as=0.4026p ps=2.71u w=0.915u l=0.5u
X1 VSS A2 a_67_756# VPW nfet_05v0 ad=0.3828p pd=2.08u as=0.1716p ps=1.18u w=0.66u l=0.6u
X2 VDD A2 a_255_756# VNW pfet_05v0 ad=0.57645p pd=2.69u as=0.2379p ps=1.435u w=0.915u l=0.5u
X3 Z a_67_756# VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.3828p ps=2.08u w=1.32u l=0.6u
X4 Z a_67_756# VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.57645p ps=2.69u w=1.83u l=0.5u
X5 a_67_756# A1 VSS VPW nfet_05v0 ad=0.1716p pd=1.18u as=0.2904p ps=2.2u w=0.66u l=0.6u
.ends

.subckt Register_unitcell$2 VDDd out q default d phi2 en phi1 VSSd
XDFF_2phase_1$3_0 VDDd d q phi1 phi2 VSSd DFF_2phase_1$3
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$3_0 en VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1$3_0/ZN
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1$3
Xgf180mcu_fd_sc_mcu9t5v0__and2_1$3_0 gf180mcu_fd_sc_mcu9t5v0__inv_1$3_0/ZN default
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1$3_0/A1 VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1$3
Xgf180mcu_fd_sc_mcu9t5v0__and2_1$3_1 q en VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1$3_0/A2
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1$3
Xgf180mcu_fd_sc_mcu9t5v0__or2_1$3_0 gf180mcu_fd_sc_mcu9t5v0__or2_1$3_0/A1 gf180mcu_fd_sc_mcu9t5v0__or2_1$3_0/A2
+ VDDd VSSd out VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1$3
.ends

.subckt SRegister_10$1 out[1] out[2] out[3] out[8] d q default10 default9 default8
+ default7 default6 default5 default4 default3 default2 default1 out[9] out[6] out[4]
+ out[10] out[7] en phi2 phi1 out[5] VDDd VSSd
XRegister_unitcell$2_0 VDDd out[2] Register_unitcell$2_7/d default2 Register_unitcell$2_6/q
+ phi2 en phi1 VSSd Register_unitcell$2
XRegister_unitcell$2_1 VDDd out[6] Register_unitcell$2_2/d default6 Register_unitcell$2_9/q
+ phi2 en phi1 VSSd Register_unitcell$2
XRegister_unitcell$2_3 VDDd out[8] Register_unitcell$2_4/d default8 Register_unitcell$2_3/d
+ phi2 en phi1 VSSd Register_unitcell$2
XRegister_unitcell$2_2 VDDd out[7] Register_unitcell$2_3/d default7 Register_unitcell$2_2/d
+ phi2 en phi1 VSSd Register_unitcell$2
XRegister_unitcell$2_4 VDDd out[9] Register_unitcell$2_5/d default9 Register_unitcell$2_4/d
+ phi2 en phi1 VSSd Register_unitcell$2
XRegister_unitcell$2_5 VDDd out[10] q default10 Register_unitcell$2_5/d phi2 en phi1
+ VSSd Register_unitcell$2
XRegister_unitcell$2_6 VDDd out[1] Register_unitcell$2_6/q default1 d phi2 en phi1
+ VSSd Register_unitcell$2
XRegister_unitcell$2_7 VDDd out[3] Register_unitcell$2_8/d default3 Register_unitcell$2_7/d
+ phi2 en phi1 VSSd Register_unitcell$2
XRegister_unitcell$2_8 VDDd out[4] Register_unitcell$2_9/d default4 Register_unitcell$2_8/d
+ phi2 en phi1 VSSd Register_unitcell$2
XRegister_unitcell$2_9 VDDd out[5] Register_unitcell$2_9/q default5 Register_unitcell$2_9/d
+ phi2 en phi1 VSSd Register_unitcell$2
.ends

.subckt pfet$315 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$337 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$335 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$333 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$318 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$316 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$314 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$336 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$334 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$317 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt asc_hysteresis_buffer$5 vss in vdd out
Xpfet$315_0 vdd vdd m1_884_42# m1_348_648# pfet$315
Xnfet$337_0 m1_1156_42# vss m1_884_42# vss nfet$337
Xnfet$335_0 in vss m1_348_648# vss nfet$335
Xnfet$333_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$333
Xpfet$318_0 vdd vdd m1_884_42# m1_1156_42# pfet$318
Xpfet$316_0 vdd vdd m1_348_648# in pfet$316
Xpfet$314_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd
+ m1_884_42# m1_884_42# pfet$314
Xnfet$336_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$336
Xnfet$334_0 m1_348_648# vss m1_884_42# vss nfet$334
Xpfet$317_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$317
.ends

.subckt pfet$320 a_28_460# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_460# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt nfet$339 a_30_n132# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt nfet$338 a_n84_0# a_94_0# a_30_460# VSUBS
X0 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$319 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=2.6p pd=9.3u as=2.6p ps=9.3u w=4u l=0.28u
.ends

.subckt SCHMITT$2 VDD VSS IN OUT
Xpfet$320_0 OUT VDD m1_596_1544# VSS pfet$320
Xnfet$339_0 OUT m1_592_402# VDD VSS nfet$339
Xnfet$338_0 m1_592_402# OUT IN VSS nfet$338
Xnfet$338_1 VSS m1_592_402# IN VSS nfet$338
Xpfet$319_1 IN VDD VDD m1_596_1544# pfet$319
Xpfet$319_0 IN VDD m1_596_1544# OUT pfet$319
.ends

.subckt scan_chain ENd CLKd out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8]
+ out[9] out[10] out[20] out[19] out[18] out[17] out[16] out[15] out[14] out[13] out[12]
+ out[11] out[21] out[22] out[23] out[24] out[25] out[26] out[27] out[28] out[29]
+ out[30] out[40] out[39] out[38] out[37] out[36] out[35] out[34] out[33] out[32]
+ out[31] out[41] out[42] out[43] out[44] out[45] out[46] out[47] out[48] out[49]
+ out[50] DATAd VDDd VSSd
Xqw_NOLclk$1_0 SCHMITT$2_0/OUT VDDd VSSd qw_NOLclk$1_0/PHI_1 qw_NOLclk$1_0/PHI_2 qw_NOLclk$1
XSRegister_10$1_0 out[31] out[32] out[33] out[38] SRegister_10$1_3/q SRegister_10$1_2/d
+ VSSd VSSd VDDd VSSd VSSd VDDd VDDd VSSd VSSd VSSd out[39] out[36] out[34] out[40]
+ out[37] SRegister_10$1_4/en qw_NOLclk$1_0/PHI_2 qw_NOLclk$1_0/PHI_1 out[35] VDDd
+ VSSd SRegister_10$1
XSRegister_10$1_1 out[11] out[12] out[13] out[18] SRegister_10$1_4/q SRegister_10$1_3/d
+ VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd out[19] out[16] out[14] out[20]
+ out[17] SRegister_10$1_4/en qw_NOLclk$1_0/PHI_2 qw_NOLclk$1_0/PHI_1 out[15] VDDd
+ VSSd SRegister_10$1
XSRegister_10$1_2 out[41] out[42] out[43] out[48] SRegister_10$1_2/d SRegister_10$1_2/q
+ VSSd VSSd VSSd VSSd VDDd VSSd VSSd VDDd VDDd VSSd out[49] out[46] out[44] out[50]
+ out[47] SRegister_10$1_4/en qw_NOLclk$1_0/PHI_2 qw_NOLclk$1_0/PHI_1 out[45] VDDd
+ VSSd SRegister_10$1
XSRegister_10$1_3 out[21] out[22] out[23] out[28] SRegister_10$1_3/d SRegister_10$1_3/q
+ VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd out[29] out[26] out[24] out[30]
+ out[27] SRegister_10$1_4/en qw_NOLclk$1_0/PHI_2 qw_NOLclk$1_0/PHI_1 out[25] VDDd
+ VSSd SRegister_10$1
XSRegister_10$1_4 out[1] out[2] out[3] out[8] SRegister_10$1_4/d SRegister_10$1_4/q
+ VSSd VSSd VSSd VSSd VDDd VSSd VSSd VSSd VSSd VSSd out[9] out[6] out[4] out[10] out[7]
+ SRegister_10$1_4/en qw_NOLclk$1_0/PHI_2 qw_NOLclk$1_0/PHI_1 out[5] VDDd VSSd SRegister_10$1
Xasc_hysteresis_buffer$5_0 VSSd CLKd VDDd SCHMITT$2_0/IN asc_hysteresis_buffer$5
XSCHMITT$2_0 VDDd VSSd SCHMITT$2_0/IN SCHMITT$2_0/OUT SCHMITT$2
Xasc_hysteresis_buffer$5_1 VSSd ENd VDDd SRegister_10$1_4/en asc_hysteresis_buffer$5
Xasc_hysteresis_buffer$5_2 VSSd DATAd VDDd SRegister_10$1_4/d asc_hysteresis_buffer$5
.ends

.subckt pfet$345 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$343 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$367 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$365 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$346 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$344 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$368 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$366 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$364 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$347 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt asc_hysteresis_buffer$6 vss in vdd out
Xpfet$345_0 vdd vdd m1_348_648# in pfet$345
Xpfet$343_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd
+ m1_884_42# m1_884_42# pfet$343
Xnfet$367_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$367
Xnfet$365_0 m1_348_648# vss m1_884_42# vss nfet$365
Xpfet$346_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$346
Xpfet$344_0 vdd vdd m1_884_42# m1_348_648# pfet$344
Xnfet$368_0 m1_1156_42# vss m1_884_42# vss nfet$368
Xnfet$366_0 in vss m1_348_648# vss nfet$366
Xnfet$364_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$364
Xpfet$347_0 vdd vdd m1_884_42# m1_1156_42# pfet$347
.ends

.subckt top_level_20250919_sc en clk data ext_pfd_div ext_pfd_ref ext_pfd_down ext_pfd_up
+ i_cp_100u filter_in filter_out ext_vco_in div_in ext_vco_out up out down lock ref
+ div_out div_def VDDd VSSd
Xtop_level_20250912_nosc_0 i_cp_100u asc_hysteresis_buffer$6_0/out scan_chain_0/out[42]
+ scan_chain_0/out[43] scan_chain_0/out[44] scan_chain_0/out[45] scan_chain_0/out[46]
+ scan_chain_0/out[47] scan_chain_0/out[48] scan_chain_0/out[49] scan_chain_0/out[50]
+ div_out div_in scan_chain_0/out[41] scan_chain_0/out[40] scan_chain_0/out[39] scan_chain_0/out[38]
+ scan_chain_0/out[37] scan_chain_0/out[36] scan_chain_0/out[35] scan_chain_0/out[34]
+ scan_chain_0/out[33] lock ref ext_pfd_div ext_pfd_ref ext_pfd_up ext_pfd_down scan_chain_0/out[1]
+ scan_chain_0/out[2] down scan_chain_0/out[6] scan_chain_0/out[5] scan_chain_0/out[4]
+ scan_chain_0/out[3] filter_in filter_out scan_chain_0/out[32] scan_chain_0/out[31]
+ scan_chain_0/out[26] scan_chain_0/out[17] scan_chain_0/out[16] scan_chain_0/out[25]
+ scan_chain_0/out[15] scan_chain_0/out[24] scan_chain_0/out[14] scan_chain_0/out[13]
+ scan_chain_0/out[12] scan_chain_0/out[11] scan_chain_0/out[10] scan_chain_0/out[9]
+ scan_chain_0/out[23] scan_chain_0/out[22] scan_chain_0/out[21] scan_chain_0/out[20]
+ scan_chain_0/out[19] scan_chain_0/out[18] scan_chain_0/out[7] scan_chain_0/out[8]
+ VCOfinal_0/fout VCOfinal_0/irefn VCOfinal_0/vin ext_vco_out up VSSd VCOfinal_0/irefp
+ VCOfinal_0/iref200 out ext_vco_in VDDd top_level_20250912_nosc
XVCOfinal_0 VCOfinal_0/s3 VCOfinal_0/s0 VCOfinal_0/s1 VCOfinal_0/s2 VCOfinal_0/iref200
+ VCOfinal_0/fout VCOfinal_0/foutb VSSd VCOfinal_0/irefn VCOfinal_0/irefp VCOfinal_0/vin
+ VSSd VDDd VCOfinal
Xscan_chain_0 en clk scan_chain_0/out[1] scan_chain_0/out[2] scan_chain_0/out[3] scan_chain_0/out[4]
+ scan_chain_0/out[5] scan_chain_0/out[6] scan_chain_0/out[7] scan_chain_0/out[8]
+ scan_chain_0/out[9] scan_chain_0/out[10] scan_chain_0/out[20] scan_chain_0/out[19]
+ scan_chain_0/out[18] scan_chain_0/out[17] scan_chain_0/out[16] scan_chain_0/out[15]
+ scan_chain_0/out[14] scan_chain_0/out[13] scan_chain_0/out[12] scan_chain_0/out[11]
+ scan_chain_0/out[21] scan_chain_0/out[22] scan_chain_0/out[23] scan_chain_0/out[24]
+ scan_chain_0/out[25] scan_chain_0/out[26] VCOfinal_0/s0 VCOfinal_0/s1 VCOfinal_0/s2
+ VCOfinal_0/s3 scan_chain_0/out[40] scan_chain_0/out[39] scan_chain_0/out[38] scan_chain_0/out[37]
+ scan_chain_0/out[36] scan_chain_0/out[35] scan_chain_0/out[34] scan_chain_0/out[33]
+ scan_chain_0/out[32] scan_chain_0/out[31] scan_chain_0/out[41] scan_chain_0/out[42]
+ scan_chain_0/out[43] scan_chain_0/out[44] scan_chain_0/out[45] scan_chain_0/out[46]
+ scan_chain_0/out[47] scan_chain_0/out[48] scan_chain_0/out[49] scan_chain_0/out[50]
+ data VDDd VSSd scan_chain
Xasc_hysteresis_buffer$6_0 VSSd div_def VDDd asc_hysteresis_buffer$6_0/out asc_hysteresis_buffer$6
.ends

.subckt top_level_20250919_final ref ext_pfd_div ext_pfd_ref ext_pfd_up ext_pfd_down
+ lock i_cp_100u up down filter_in ext_vco_out ext_vco_in filter_out out div_in div_out
+ div_def clk data en VSSd VDDd
Xppolyf_u_resistor$6_0 VSSd top_level_20250919_sc_0/en VSSd ppolyf_u_resistor$6
XDECAP_LARGE_0 VDDd VSSd DECAP_LARGE
Xio_secondary_3p3_0 ref VDDd VSSd io_secondary_3p3_0/to_gate io_secondary_3p3
Xio_secondary_3p3_1 i_cp_100u VDDd VSSd io_secondary_3p3_1/to_gate io_secondary_3p3
Xio_secondary_3p3_2 div_def VDDd VSSd io_secondary_3p3_2/to_gate io_secondary_3p3
Xio_secondary_3p3_4 data VDDd VSSd io_secondary_3p3_4/to_gate io_secondary_3p3
Xio_secondary_3p3_3 clk VDDd VSSd io_secondary_3p3_3/to_gate io_secondary_3p3
Xio_secondary_3p3_5 en VDDd VSSd top_level_20250919_sc_0/en io_secondary_3p3
Xtop_level_20250919_sc_0 top_level_20250919_sc_0/en io_secondary_3p3_3/to_gate io_secondary_3p3_4/to_gate
+ ext_pfd_div ext_pfd_ref ext_pfd_down ext_pfd_up io_secondary_3p3_1/to_gate filter_in
+ filter_out ext_vco_in div_in ext_vco_out up out down lock io_secondary_3p3_0/to_gate
+ div_out io_secondary_3p3_2/to_gate VDDd VSSd top_level_20250919_sc
.ends

