* Extracted by KLayout with GF180MCU LVS runset on : 09/08/2025 17:31

.SUBCKT asc_NAND VSS B OUT A VDD
M$1 VDD B OUT VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$2 OUT A VDD VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$3 \$2 B VSS VSS nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U PD=4.74U
M$5 \$2 A OUT VSS nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U PD=4.74U
.ENDS asc_NAND
