* Extracted by KLayout with GF180MCU LVS runset on : 09/08/2025 17:36

.SUBCKT asc_NOR VSS OUT A B VDD
M$1 \$9 A VDD VDD pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U PD=10.82U
M$3 \$9 B OUT VDD pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U PD=10.82U
M$5 VSS A OUT VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$6 OUT B VSS VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
.ENDS asc_NOR
