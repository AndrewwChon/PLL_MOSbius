* Extracted by KLayout with GF180MCU LVS runset on : 15/09/2025 00:21

.SUBCKT asc_dual_psd_def_20250809 sd9 sd8 sd7 sd6 sd5 sd4 sd3 sd2 sd1 vss fout
+ define fin pd1 pd2 pd3 pd4 pd5 pd6 pd7 pd8 pd9
M$1 \$544 sd9 \$76 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$2 \$544 \$119 \$77 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$3 \$77 \$120 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$4 \$78 \$2 \$120 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$5 \$544 \$121 \$78 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$6 \$80 \$79 \$121 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$7 \$544 \$77 \$80 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$8 \$544 \$2 \$79 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$9 \$544 sd8 \$3 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$10 \$544 \$447 \$81 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$11 \$81 \$123 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$12 \$82 \$4 \$123 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$13 \$544 \$124 \$82 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$14 \$84 \$83 \$124 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$15 \$544 \$81 \$84 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$16 \$544 \$4 \$83 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$17 \$544 sd7 \$85 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$18 \$544 \$126 \$86 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$19 \$86 \$127 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$20 \$87 \$5 \$127 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$21 \$544 \$128 \$87 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$22 \$89 \$88 \$128 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$23 \$544 \$86 \$89 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$24 \$544 \$5 \$88 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$25 \$544 sd6 \$90 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$26 \$544 \$130 \$91 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$27 \$91 \$131 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$28 \$92 \$6 \$131 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$29 \$544 \$132 \$92 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$30 \$94 \$93 \$132 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$31 \$544 \$91 \$94 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$32 \$544 \$6 \$93 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$33 \$544 sd5 \$7 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$34 \$544 \$135 \$134 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$35 \$134 \$136 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$36 \$95 \$8 \$136 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$37 \$544 \$137 \$95 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$38 \$97 \$96 \$137 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$39 \$544 \$134 \$97 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$40 \$544 \$8 \$96 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$41 \$544 sd4 \$98 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$42 \$544 \$139 \$99 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$43 \$99 \$140 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$44 \$100 \$9 \$140 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$45 \$544 \$141 \$100 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$46 \$102 \$101 \$141 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$47 \$544 \$99 \$102 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$48 \$544 \$9 \$101 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$49 \$544 sd3 \$103 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$50 \$544 \$143 \$104 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$51 \$104 \$144 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$52 \$105 \$10 \$144 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$53 \$544 \$145 \$105 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$54 \$107 \$106 \$145 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$55 \$544 \$104 \$107 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$56 \$544 \$10 \$106 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$57 \$544 sd2 \$108 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$58 \$544 \$466 \$109 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$59 \$109 \$147 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$60 \$110 \$11 \$147 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$61 \$544 \$148 \$110 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$62 \$112 \$111 \$148 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$63 \$544 \$109 \$112 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$64 \$544 \$11 \$111 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$65 \$544 sd1 \$113 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$66 \$544 \$150 \$114 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$67 \$114 \$151 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$68 \$115 \$12 \$151 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$69 \$544 \$152 \$115 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$70 \$117 \$116 \$152 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$71 \$544 \$114 \$117 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$72 \$544 \$12 \$116 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$73 \$544 \$77 \$442 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$74 \$443 \$77 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$75 \$120 \$79 \$443 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$76 \$119 \$1 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$77 \$544 \$119 \$444 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$78 \$444 \$78 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$79 \$121 \$2 \$444 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$80 \$544 \$445 \$2 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$81 \$544 \$81 \$445 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$82 \$446 \$81 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$83 \$123 \$83 \$446 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$84 \$447 \$1 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$85 \$544 \$447 \$448 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$86 \$448 \$82 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$87 \$124 \$4 \$448 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$88 \$544 \$449 \$4 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$89 \$544 \$86 \$449 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$90 \$450 \$86 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$91 \$127 \$88 \$450 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$92 \$126 \$1 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$93 \$544 \$126 \$451 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$94 \$451 \$87 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$95 \$128 \$5 \$451 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$96 \$544 \$452 \$5 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$97 \$544 \$91 \$452 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$98 \$453 \$91 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$99 \$131 \$93 \$453 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$100 \$130 \$1 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$101 \$544 \$130 \$454 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$102 \$454 \$92 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$103 \$132 \$6 \$454 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$104 \$544 \$455 \$6 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$105 \$544 \$134 \$455 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$106 \$456 \$134 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$107 \$136 \$96 \$456 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$108 \$135 \$1 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$109 \$544 \$135 \$457 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$110 \$457 \$95 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$111 \$137 \$8 \$457 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$112 \$544 \$458 \$8 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$113 \$544 \$99 \$458 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$114 \$459 \$99 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$115 \$140 \$101 \$459 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$116 \$139 \$1 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$117 \$544 \$139 \$460 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$118 \$460 \$100 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$119 \$141 \$9 \$460 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$120 \$544 \$461 \$9 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$121 \$544 \$104 \$461 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$122 \$462 \$104 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$123 \$144 \$106 \$462 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$124 \$143 \$1 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$125 \$544 \$143 \$463 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$126 \$463 \$105 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$127 \$145 \$10 \$463 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$128 \$544 \$464 \$10 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$129 \$544 \$109 \$464 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$130 \$465 \$109 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$131 \$147 \$111 \$465 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$132 \$466 \$1 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$133 \$544 \$466 \$467 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$134 \$467 \$110 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$135 \$148 \$11 \$467 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$136 \$544 \$468 \$11 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$137 \$544 \$114 \$468 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$138 \$469 \$114 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$139 \$151 \$116 \$469 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$140 \$150 \$1 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$141 \$544 \$150 \$470 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$142 \$470 \$115 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$143 \$152 \$12 \$470 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$144 \$544 \$471 \$12 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$145 \$738 \$787 \$737 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$147 \$738 \$1 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$149 \$544 \$740 \$739 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$150 \$544 \$788 \$740 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$151 \$740 \$680 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$152 \$742 \$744 \$741 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$154 \$742 \$743 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$156 \$544 \$688 \$743 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$157 \$743 \$687 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$158 \$544 \$686 \$744 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$159 \$744 \$685 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$160 \$745 \$442 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$161 \$746 \$745 \$680 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$163 \$747 \$442 \$680 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$165 \$747 \$76 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$167 \$746 \$748 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$169 \$544 \$76 \$748 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$170 \$749 \$445 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$171 \$750 \$749 \$681 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$173 \$751 \$445 \$681 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$175 \$751 \$3 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$177 \$750 \$752 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$179 \$544 \$3 \$752 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$180 \$753 \$449 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$181 \$754 \$753 \$682 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$183 \$755 \$449 \$682 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$185 \$755 \$85 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$187 \$754 \$756 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$189 \$544 \$85 \$756 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$190 \$757 \$452 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$191 \$758 \$757 \$683 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$193 \$759 \$452 \$683 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$195 \$759 \$90 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$197 \$758 \$760 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$199 \$544 \$90 \$760 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$200 \$761 \$455 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$201 \$762 \$761 \$684 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$203 \$763 \$455 \$684 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$205 \$763 \$7 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$207 \$762 \$764 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$209 \$544 \$7 \$764 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$210 \$765 \$458 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$211 \$766 \$765 \$685 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$213 \$767 \$458 \$685 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$215 \$767 \$98 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$217 \$766 \$768 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$219 \$544 \$98 \$768 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$220 \$769 \$461 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$221 \$770 \$769 \$686 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$223 \$771 \$461 \$686 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$225 \$771 \$103 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$227 \$770 \$772 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$229 \$544 \$103 \$772 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$230 \$773 \$464 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$231 \$774 \$773 \$687 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$233 \$775 \$464 \$687 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$235 \$775 \$108 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$237 \$774 \$776 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$239 \$544 \$108 \$776 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$240 \$777 \$468 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$241 \$778 \$777 \$688 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$243 \$779 \$468 \$688 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$245 \$779 \$113 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$247 \$778 \$780 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$249 \$544 \$113 \$780 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$250 \$544 \$1081 \$781 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$251 \$781 \$1079 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$252 \$544 \$1077 \$782 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$253 \$782 \$1075 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$254 \$783 \$782 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$256 \$783 \$781 \$784 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$258 \$544 \$784 \$785 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$259 \$785 \$865 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$260 \$786 \$785 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$261 \$544 \$789 \$1 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$262 \$1217 \$739 \$787 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$264 \$1217 \$737 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$266 \$544 \$1088 \$788 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$267 \$544 \$741 \$1088 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$268 \$1088 \$1089 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$269 \$1218 \$1064 \$1089 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$271 \$1218 \$1090 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$273 \$544 \$684 \$1090 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$274 \$1090 \$683 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$275 \$544 \$682 \$1064 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$276 \$1064 \$681 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$277 \$1092 \$1091 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$278 \$1219 \$1092 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$280 \$1220 \$1091 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$282 \$1220 \$1094 \$1067 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$284 \$1219 \$1095 \$1067 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$286 \$544 \$1094 \$1095 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$287 \$1097 \$1096 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$288 \$1221 \$1097 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$290 \$1222 \$1096 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$292 \$1222 \$1099 \$1069 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$294 \$1221 \$1100 \$1069 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$296 \$544 \$1099 \$1100 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$297 \$1102 \$1101 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$298 \$1223 \$1102 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$300 \$1224 \$1101 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$302 \$1224 \$1104 \$1071 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$304 \$1223 \$1105 \$1071 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$306 \$544 \$1104 \$1105 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$307 \$1107 \$1106 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$308 \$1225 \$1107 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$310 \$1226 \$1106 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$312 \$1226 \$1109 \$1073 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$314 \$1225 \$1110 \$1073 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$316 \$544 \$1109 \$1110 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$317 \$1112 \$1111 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$318 \$1227 \$1112 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$320 \$1228 \$1111 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$322 \$1228 \$1114 \$1075 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$324 \$1227 \$1115 \$1075 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$326 \$544 \$1114 \$1115 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$327 \$1117 \$1116 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$328 \$1229 \$1117 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$330 \$1230 \$1116 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$332 \$1230 \$1119 \$1077 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$334 \$1229 \$1120 \$1077 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$336 \$544 \$1119 \$1120 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$337 \$1122 \$1121 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$338 \$1231 \$1122 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$340 \$1232 \$1121 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$342 \$1232 \$1124 \$1079 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$344 \$1231 \$1125 \$1079 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$346 \$544 \$1124 \$1125 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$347 \$1127 \$1126 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$348 \$1233 \$1127 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$350 \$1234 \$1126 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$352 \$1234 \$1129 \$1081 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$354 \$1233 \$1130 \$1081 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$356 \$544 \$1129 \$1130 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$357 \$1132 \$1131 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$358 \$1235 \$1132 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$360 \$1236 \$1131 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$362 \$1236 \$1134 \$1083 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$364 \$1235 \$1135 \$1083 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$366 \$544 \$1134 \$1135 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$367 \$544 \$1073 \$1136 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$368 \$1136 \$1071 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$369 \$544 \$1069 \$1137 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$370 \$1137 \$1067 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$371 \$1237 \$1137 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$373 \$1237 \$1136 \$865 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$375 \$544 \$1083 \$1138 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$376 \$1138 \$786 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$377 fout \$1138 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$378 \$1238 fout \$789 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$380 \$1238 define \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$382 \$1624 \$1442 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$383 \$1442 fin \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$384 \$1904 \$471 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$385 \$1444 \$1442 \$1443 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$386 \$1443 \$1624 \$1904 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$387 \$544 \$1509 \$1444 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$388 \$1509 \$1443 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$389 \$1444 \$1445 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$390 \$1446 \$1442 \$1509 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$391 \$544 vss \$1445 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$392 \$544 \$1446 \$1510 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$393 \$1447 \$1624 \$1446 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$394 \$544 \$1510 \$1447 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$395 \$1510 \$1445 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$396 \$1448 \$1510 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$397 \$544 \$1905 \$1514 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$398 \$544 \$471 \$1905 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$399 \$1449 \$1448 \$544 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$401 \$1449 \$737 \$1450 \$544 pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$403 \$1905 \$1451 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$404 \$1451 \$1450 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$405 \$544 \$471 \$1906 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$406 \$544 \$1511 \$471 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$407 \$1907 \$471 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$408 \$1512 \$1636 \$1907 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$409 \$471 \$1512 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$410 \$1511 vss \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$411 \$1452 \$1363 \$1512 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$412 \$544 \$1511 \$1908 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$413 \$544 \$1513 \$1452 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$414 \$1453 \$1636 \$1513 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$415 \$1908 \$1452 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$416 \$1513 \$1363 \$1908 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$417 \$544 \$1514 \$1453 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$418 \$544 fin \$1363 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$419 \$544 \$1363 \$1636 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$420 \$1625 \$1454 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$421 \$1454 \$471 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$422 \$1909 \$1516 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$423 \$1456 \$1454 \$1455 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$424 \$544 \$1515 \$1456 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$425 \$1455 \$1625 \$1909 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$426 \$1515 \$1455 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$427 \$1456 \$1457 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$428 \$1458 \$1454 \$1515 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$429 \$544 \$1 \$1457 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$430 \$544 \$1458 \$1516 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$431 \$1459 \$1625 \$1458 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$432 \$544 \$1516 \$1459 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$433 \$1516 \$1457 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$434 \$1091 pd1 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$435 \$1094 \$1516 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$436 \$1626 \$1460 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$437 \$1460 \$1094 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$438 \$1910 \$1518 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$439 \$1462 \$1460 \$1461 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$440 \$1461 \$1626 \$1910 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$441 \$544 \$1517 \$1462 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$442 \$1517 \$1461 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$443 \$1462 \$1463 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$444 \$1464 \$1460 \$1517 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$445 \$544 \$1 \$1463 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$446 \$544 \$1464 \$1518 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$447 \$1465 \$1626 \$1464 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$448 \$544 \$1518 \$1465 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$449 \$1518 \$1463 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$450 \$1099 \$1518 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$451 \$1096 pd2 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$452 \$1627 \$1466 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$453 \$1466 \$1099 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$454 \$1911 \$1520 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$455 \$1468 \$1466 \$1467 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$456 \$1467 \$1627 \$1911 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$457 \$544 \$1519 \$1468 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$458 \$1519 \$1467 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$459 \$1468 \$1469 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$460 \$1470 \$1466 \$1519 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$461 \$544 \$1 \$1469 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$462 \$544 \$1470 \$1520 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$463 \$1471 \$1627 \$1470 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$464 \$544 \$1520 \$1471 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$465 \$1520 \$1469 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$466 \$1104 \$1520 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$467 \$1101 pd3 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$468 \$1628 \$1472 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$469 \$1472 \$1104 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$470 \$1912 \$1522 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$471 \$1474 \$1472 \$1473 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$472 \$1473 \$1628 \$1912 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$473 \$544 \$1521 \$1474 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$474 \$1521 \$1473 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$475 \$1474 \$1475 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$476 \$1476 \$1472 \$1521 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$477 \$544 \$1 \$1475 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$478 \$544 \$1476 \$1522 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$479 \$1477 \$1628 \$1476 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$480 \$544 \$1522 \$1477 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$481 \$1522 \$1475 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$482 \$1106 pd4 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$483 \$1109 \$1522 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$484 \$1629 \$1478 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$485 \$1478 \$1109 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$486 \$1913 \$1524 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$487 \$1480 \$1478 \$1479 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$488 \$544 \$1523 \$1480 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$489 \$1479 \$1629 \$1913 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$490 \$1523 \$1479 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$491 \$1480 \$1481 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$492 \$1482 \$1478 \$1523 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$493 \$544 \$1 \$1481 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$494 \$544 \$1482 \$1524 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$495 \$1483 \$1629 \$1482 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$496 \$544 \$1524 \$1483 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$497 \$1524 \$1481 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$498 \$1114 \$1524 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$499 \$1111 pd5 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$500 \$1630 \$1484 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$501 \$1484 \$1114 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$502 \$1914 \$1526 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$503 \$1486 \$1484 \$1485 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$504 \$544 \$1525 \$1486 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$505 \$1485 \$1630 \$1914 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$506 \$1525 \$1485 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$507 \$1486 \$1487 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$508 \$1488 \$1484 \$1525 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$509 \$544 \$1 \$1487 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$510 \$544 \$1488 \$1526 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$511 \$1489 \$1630 \$1488 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$512 \$544 \$1526 \$1489 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$513 \$1526 \$1487 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$514 \$1116 pd6 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$515 \$1119 \$1526 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$516 \$1631 \$1490 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$517 \$1490 \$1119 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$518 \$1915 \$1528 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$519 \$1492 \$1490 \$1491 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$520 \$544 \$1527 \$1492 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$521 \$1491 \$1631 \$1915 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$522 \$1527 \$1491 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$523 \$1492 \$1493 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$524 \$1494 \$1490 \$1527 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$525 \$544 \$1 \$1493 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$526 \$544 \$1494 \$1528 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$527 \$1495 \$1631 \$1494 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$528 \$544 \$1528 \$1495 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$529 \$1528 \$1493 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$530 \$1121 pd7 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$531 \$1124 \$1528 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$532 \$1632 \$1496 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$533 \$1496 \$1124 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$534 \$1916 \$1530 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$535 \$1498 \$1496 \$1497 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$536 \$544 \$1529 \$1498 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$537 \$1497 \$1632 \$1916 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$538 \$1529 \$1497 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$539 \$1498 \$1499 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$540 \$1500 \$1496 \$1529 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$541 \$544 \$1 \$1499 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$542 \$544 \$1500 \$1530 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$543 \$1501 \$1632 \$1500 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$544 \$544 \$1530 \$1501 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$545 \$1530 \$1499 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$546 \$1129 \$1530 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$547 \$1126 pd8 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$548 \$1633 \$1502 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$549 \$1502 \$1129 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$550 \$1917 \$1532 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$551 \$1504 \$1502 \$1503 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$552 \$544 \$1531 \$1504 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$553 \$1503 \$1633 \$1917 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$554 \$1531 \$1503 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$555 \$1504 \$1505 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$556 \$1506 \$1502 \$1531 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$557 \$544 \$1 \$1505 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$558 \$544 \$1506 \$1532 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$559 \$1507 \$1633 \$1506 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$560 \$544 \$1532 \$1507 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$561 \$1532 \$1505 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$562 \$1134 \$1532 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$563 \$1131 pd9 \$544 \$544 pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$564 vss sd9 \$76 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$565 \$226 \$119 \$77 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$567 \$226 \$120 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$569 \$78 \$79 \$120 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$570 vss \$121 \$78 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$571 \$80 \$2 \$121 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$572 vss \$77 \$80 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$573 vss \$2 \$79 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$574 vss sd8 \$3 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$575 \$227 \$447 \$81 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$577 \$227 \$123 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$579 \$82 \$83 \$123 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$580 vss \$124 \$82 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$581 \$84 \$4 \$124 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$582 vss \$81 \$84 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$583 vss \$4 \$83 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$584 vss sd7 \$85 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$585 \$228 \$126 \$86 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$587 \$228 \$127 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$589 \$87 \$88 \$127 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$590 vss \$128 \$87 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$591 \$89 \$5 \$128 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$592 vss \$86 \$89 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$593 vss \$5 \$88 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$594 vss sd6 \$90 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$595 \$229 \$130 \$91 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$597 \$229 \$131 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$599 \$92 \$93 \$131 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$600 vss \$132 \$92 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$601 \$94 \$6 \$132 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$602 vss \$91 \$94 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$603 vss \$6 \$93 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$604 vss sd5 \$7 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$605 \$230 \$135 \$134 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$607 \$230 \$136 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$609 \$95 \$96 \$136 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$610 vss \$137 \$95 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$611 \$97 \$8 \$137 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$612 vss \$134 \$97 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$613 vss \$8 \$96 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$614 vss sd4 \$98 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$615 \$231 \$139 \$99 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$617 \$231 \$140 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$619 \$100 \$101 \$140 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$620 vss \$141 \$100 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$621 \$102 \$9 \$141 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$622 vss \$99 \$102 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$623 vss \$9 \$101 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$624 vss sd3 \$103 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$625 \$232 \$143 \$104 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$627 \$232 \$144 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$629 \$105 \$106 \$144 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$630 vss \$145 \$105 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$631 \$107 \$10 \$145 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$632 vss \$104 \$107 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$633 vss \$10 \$106 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$634 vss sd2 \$108 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$635 \$233 \$466 \$109 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$637 \$233 \$147 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$639 \$110 \$111 \$147 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$640 vss \$148 \$110 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$641 \$112 \$11 \$148 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$642 vss \$109 \$112 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$643 vss \$11 \$111 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$644 vss sd1 \$113 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$645 \$234 \$150 \$114 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$647 \$234 \$151 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$649 \$115 \$116 \$151 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$650 vss \$152 \$115 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$651 \$117 \$12 \$152 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$652 vss \$114 \$117 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$653 vss \$12 \$116 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$654 vss \$77 \$442 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$655 \$443 \$77 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$656 \$120 \$2 \$443 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$657 \$119 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$658 \$370 \$119 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$660 \$370 \$78 \$444 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$662 \$121 \$79 \$444 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$663 vss \$445 \$2 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$664 vss \$81 \$445 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$665 \$446 \$81 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$666 \$123 \$4 \$446 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$667 \$447 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$668 \$371 \$447 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$670 \$371 \$82 \$448 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$672 \$124 \$83 \$448 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$673 vss \$449 \$4 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$674 vss \$86 \$449 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$675 \$450 \$86 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$676 \$127 \$5 \$450 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$677 \$126 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$678 \$372 \$126 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$680 \$372 \$87 \$451 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$682 \$128 \$88 \$451 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$683 vss \$452 \$5 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$684 vss \$91 \$452 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$685 \$453 \$91 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$686 \$131 \$6 \$453 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$687 \$130 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$688 \$373 \$130 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$690 \$373 \$92 \$454 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$692 \$132 \$93 \$454 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$693 vss \$455 \$6 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$694 vss \$134 \$455 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$695 \$456 \$134 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$696 \$136 \$8 \$456 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$697 \$135 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$698 \$374 \$135 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$700 \$374 \$95 \$457 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$702 \$137 \$96 \$457 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$703 vss \$458 \$8 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$704 vss \$99 \$458 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$705 \$459 \$99 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$706 \$140 \$9 \$459 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$707 \$139 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$708 \$375 \$139 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$710 \$375 \$100 \$460 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$712 \$141 \$101 \$460 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$713 vss \$461 \$9 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$714 vss \$104 \$461 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$715 \$462 \$104 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$716 \$144 \$10 \$462 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$717 \$143 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$718 \$376 \$143 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$720 \$376 \$105 \$463 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$722 \$145 \$106 \$463 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$723 vss \$464 \$10 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$724 vss \$109 \$464 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$725 \$465 \$109 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$726 \$147 \$11 \$465 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$727 \$466 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$728 \$377 \$466 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$730 \$377 \$110 \$467 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$732 \$148 \$111 \$467 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$733 vss \$468 \$11 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$734 vss \$114 \$468 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$735 \$469 \$114 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$736 \$151 \$12 \$469 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$737 \$150 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$738 \$378 \$150 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$740 \$378 \$115 \$470 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$742 \$152 \$116 \$470 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$743 vss \$471 \$12 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$744 vss \$787 \$737 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$745 \$737 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$746 vss \$740 \$739 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$747 \$868 \$788 \$740 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$749 \$868 \$680 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$751 vss \$744 \$741 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$752 \$741 \$743 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$753 \$869 \$688 \$743 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$755 \$869 \$687 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$757 \$870 \$686 \$744 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$759 \$870 \$685 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$761 \$745 \$442 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$762 \$871 \$745 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$764 \$872 \$442 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$766 \$871 \$76 \$680 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$768 \$872 \$748 \$680 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$770 vss \$76 \$748 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$771 \$749 \$445 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$772 \$873 \$749 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$774 \$874 \$445 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$776 \$873 \$3 \$681 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$778 \$874 \$752 \$681 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$780 vss \$3 \$752 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$781 \$753 \$449 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$782 \$875 \$753 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$784 \$876 \$449 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$786 \$875 \$85 \$682 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$788 \$876 \$756 \$682 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$790 vss \$85 \$756 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$791 \$757 \$452 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$792 \$877 \$757 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$794 \$878 \$452 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$796 \$877 \$90 \$683 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$798 \$878 \$760 \$683 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$800 vss \$90 \$760 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$801 \$761 \$455 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$802 \$879 \$761 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$804 \$880 \$455 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$806 \$879 \$7 \$684 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$808 \$880 \$764 \$684 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$810 vss \$7 \$764 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$811 \$765 \$458 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$812 \$881 \$765 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$814 \$882 \$458 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$816 \$881 \$98 \$685 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$818 \$882 \$768 \$685 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$820 vss \$98 \$768 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$821 \$769 \$461 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$822 \$883 \$769 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$824 \$884 \$461 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$826 \$883 \$103 \$686 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$828 \$884 \$772 \$686 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$830 vss \$103 \$772 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$831 \$773 \$464 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$832 \$885 \$773 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$834 \$886 \$464 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$836 \$885 \$108 \$687 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$838 \$886 \$776 \$687 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$840 vss \$108 \$776 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$841 \$777 \$468 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$842 \$887 \$777 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$844 \$888 \$468 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$846 \$887 \$113 \$688 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$848 \$888 \$780 \$688 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$850 vss \$113 \$780 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$851 \$889 \$1081 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$853 \$889 \$1079 \$781 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$855 \$890 \$1077 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$857 \$890 \$1075 \$782 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$859 vss \$782 \$784 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$860 \$784 \$781 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$861 \$891 \$784 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$863 \$891 \$865 \$785 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$865 \$786 \$785 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$866 vss \$789 \$1 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$867 vss \$739 \$787 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$868 \$787 \$737 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$869 vss \$1088 \$788 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$870 \$1063 \$741 \$1088 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$872 \$1063 \$1089 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$874 vss \$1064 \$1089 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$875 \$1089 \$1090 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$876 \$1065 \$684 \$1090 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$878 \$1065 \$683 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$880 \$1066 \$682 \$1064 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$882 \$1066 \$681 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$884 \$1092 \$1091 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$885 \$1068 \$1092 \$1067 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$887 \$1093 \$1091 \$1067 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$889 \$1068 \$1094 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$891 \$1093 \$1095 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$893 vss \$1094 \$1095 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$894 \$1097 \$1096 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$895 \$1070 \$1097 \$1069 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$897 \$1098 \$1096 \$1069 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$899 \$1070 \$1099 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$901 \$1098 \$1100 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$903 vss \$1099 \$1100 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$904 \$1102 \$1101 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$905 \$1072 \$1102 \$1071 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$907 \$1103 \$1101 \$1071 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$909 \$1072 \$1104 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$911 \$1103 \$1105 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$913 vss \$1104 \$1105 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$914 \$1107 \$1106 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$915 \$1074 \$1107 \$1073 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$917 \$1108 \$1106 \$1073 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$919 \$1074 \$1109 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$921 \$1108 \$1110 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$923 vss \$1109 \$1110 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$924 \$1112 \$1111 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$925 \$1076 \$1112 \$1075 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$927 \$1113 \$1111 \$1075 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$929 \$1076 \$1114 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$931 \$1113 \$1115 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$933 vss \$1114 \$1115 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$934 \$1117 \$1116 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$935 \$1078 \$1117 \$1077 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$937 \$1118 \$1116 \$1077 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$939 \$1078 \$1119 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$941 \$1118 \$1120 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$943 vss \$1119 \$1120 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$944 \$1122 \$1121 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$945 \$1080 \$1122 \$1079 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$947 \$1123 \$1121 \$1079 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$949 \$1080 \$1124 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$951 \$1123 \$1125 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$953 vss \$1124 \$1125 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$954 \$1127 \$1126 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$955 \$1082 \$1127 \$1081 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$957 \$1128 \$1126 \$1081 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$959 \$1082 \$1129 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$961 \$1128 \$1130 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$963 vss \$1129 \$1130 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$964 \$1132 \$1131 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$965 \$1084 \$1132 \$1083 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$967 \$1133 \$1131 \$1083 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$969 \$1084 \$1134 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$971 \$1133 \$1135 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$973 vss \$1134 \$1135 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$974 \$1085 \$1073 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$976 \$1085 \$1071 \$1136 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$978 \$1086 \$1069 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$980 \$1086 \$1067 \$1137 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$982 vss \$1137 \$865 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$983 \$865 \$1136 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$984 \$1087 \$1083 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$986 \$1087 \$786 \$1138 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$988 fout \$1138 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$989 vss fout \$789 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$990 \$789 define vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$991 \$1624 \$1442 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$992 \$1442 fin vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$993 \$1904 \$471 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$994 \$1444 \$1624 \$1443 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$995 \$1443 \$1442 \$1904 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$996 \$1634 \$1509 \$1444 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$998 \$1509 \$1443 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$999 \$1634 \$1445 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1001 \$1446 \$1624 \$1509 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1002 vss vss \$1445 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1003 \$1892 \$1446 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1005 \$1447 \$1442 \$1446 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1006 \$1892 \$1445 \$1510 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1008 vss \$1510 \$1447 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1009 \$1448 \$1510 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1010 vss \$1905 \$1514 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1011 \$1893 \$471 \$1905 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1013 vss \$1448 \$1450 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1014 \$1893 \$1451 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1016 \$1450 \$737 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1017 \$1451 \$1450 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1018 vss \$471 \$1906 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1019 \$1635 \$1511 \$471 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1021 \$1907 \$471 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1022 \$1512 \$1363 \$1907 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1023 \$1635 \$1512 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1025 \$1511 vss vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1026 \$1452 \$1636 \$1512 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1027 \$1894 \$1511 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1029 vss \$1513 \$1452 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1030 \$1894 \$1452 \$1908 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1032 \$1453 \$1363 \$1513 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1033 \$1513 \$1636 \$1908 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1034 vss \$1514 \$1453 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1035 vss fin \$1363 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1036 vss \$1363 \$1636 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1037 \$1625 \$1454 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1038 \$1454 \$471 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1039 \$1909 \$1516 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1040 \$1456 \$1625 \$1455 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1041 \$1455 \$1454 \$1909 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1042 \$1637 \$1515 \$1456 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1044 \$1515 \$1455 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1045 \$1637 \$1457 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1047 \$1458 \$1625 \$1515 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1048 vss \$1 \$1457 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1049 \$1895 \$1458 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1051 \$1459 \$1454 \$1458 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1052 \$1895 \$1457 \$1516 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1054 vss \$1516 \$1459 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1055 \$1094 \$1516 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1056 \$1091 pd1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1057 \$1626 \$1460 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1058 \$1460 \$1094 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1059 \$1910 \$1518 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1060 \$1462 \$1626 \$1461 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1061 \$1638 \$1517 \$1462 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1063 \$1461 \$1460 \$1910 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1064 \$1517 \$1461 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1065 \$1638 \$1463 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1067 \$1464 \$1626 \$1517 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1068 vss \$1 \$1463 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1069 \$1896 \$1464 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1071 \$1465 \$1460 \$1464 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1072 \$1896 \$1463 \$1518 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1074 vss \$1518 \$1465 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1075 \$1099 \$1518 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1076 \$1096 pd2 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1077 \$1627 \$1466 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1078 \$1466 \$1099 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1079 \$1911 \$1520 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1080 \$1468 \$1627 \$1467 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1081 \$1467 \$1466 \$1911 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1082 \$1639 \$1519 \$1468 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1084 \$1519 \$1467 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1085 \$1639 \$1469 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1087 \$1470 \$1627 \$1519 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1088 vss \$1 \$1469 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1089 \$1897 \$1470 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1091 \$1471 \$1466 \$1470 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1092 \$1897 \$1469 \$1520 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1094 vss \$1520 \$1471 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1095 \$1104 \$1520 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1096 \$1101 pd3 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1097 \$1628 \$1472 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1098 \$1472 \$1104 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1099 \$1912 \$1522 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1100 \$1474 \$1628 \$1473 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1101 \$1473 \$1472 \$1912 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1102 \$1640 \$1521 \$1474 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1104 \$1521 \$1473 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1105 \$1640 \$1475 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1107 \$1476 \$1628 \$1521 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1108 vss \$1 \$1475 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1109 \$1898 \$1476 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1111 \$1477 \$1472 \$1476 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1112 \$1898 \$1475 \$1522 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1114 vss \$1522 \$1477 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1115 \$1109 \$1522 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1116 \$1106 pd4 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1117 \$1629 \$1478 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1118 \$1478 \$1109 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1119 \$1913 \$1524 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1120 \$1480 \$1629 \$1479 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1121 \$1641 \$1523 \$1480 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1123 \$1479 \$1478 \$1913 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1124 \$1523 \$1479 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1125 \$1641 \$1481 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1127 \$1482 \$1629 \$1523 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1128 vss \$1 \$1481 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1129 \$1899 \$1482 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1131 \$1483 \$1478 \$1482 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1132 \$1899 \$1481 \$1524 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1134 vss \$1524 \$1483 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1135 \$1114 \$1524 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1136 \$1111 pd5 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1137 \$1630 \$1484 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1138 \$1484 \$1114 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1139 \$1914 \$1526 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1140 \$1486 \$1630 \$1485 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1141 \$1485 \$1484 \$1914 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1142 \$1642 \$1525 \$1486 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1144 \$1525 \$1485 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1145 \$1642 \$1487 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1147 \$1488 \$1630 \$1525 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1148 vss \$1 \$1487 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1149 \$1900 \$1488 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1151 \$1489 \$1484 \$1488 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1152 \$1900 \$1487 \$1526 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1154 vss \$1526 \$1489 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1155 \$1119 \$1526 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1156 \$1116 pd6 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1157 \$1631 \$1490 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1158 \$1490 \$1119 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1159 \$1915 \$1528 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1160 \$1492 \$1631 \$1491 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1161 \$1643 \$1527 \$1492 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1163 \$1491 \$1490 \$1915 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1164 \$1527 \$1491 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1165 \$1643 \$1493 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1167 \$1494 \$1631 \$1527 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1168 vss \$1 \$1493 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1169 \$1901 \$1494 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1171 \$1495 \$1490 \$1494 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1172 \$1901 \$1493 \$1528 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1174 vss \$1528 \$1495 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1175 \$1124 \$1528 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1176 \$1121 pd7 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1177 \$1632 \$1496 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1178 \$1496 \$1124 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1179 \$1916 \$1530 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1180 \$1498 \$1632 \$1497 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1181 \$1644 \$1529 \$1498 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1183 \$1497 \$1496 \$1916 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1184 \$1529 \$1497 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1185 \$1644 \$1499 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1187 \$1500 \$1632 \$1529 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1188 vss \$1 \$1499 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1189 \$1902 \$1500 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1191 \$1501 \$1496 \$1500 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1192 \$1902 \$1499 \$1530 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1194 vss \$1530 \$1501 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1195 \$1126 pd8 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1196 \$1129 \$1530 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1197 \$1633 \$1502 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1198 \$1502 \$1129 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1199 \$1917 \$1532 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1200 \$1504 \$1633 \$1503 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1201 \$1645 \$1531 \$1504 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1203 \$1503 \$1502 \$1917 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1204 \$1531 \$1503 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1205 \$1645 \$1505 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1207 \$1506 \$1633 \$1531 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1208 vss \$1 \$1505 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1209 \$1903 \$1506 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1211 \$1507 \$1502 \$1506 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1212 \$1903 \$1505 \$1532 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1214 vss \$1532 \$1507 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1215 \$1131 pd9 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1216 \$1134 \$1532 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
.ENDS asc_dual_psd_def_20250809
