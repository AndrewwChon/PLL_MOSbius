** sch_path: /foss/designs/libs/secondary_esd/single_diode.sch
.subckt single_diode VDD VSS
*.PININFO VDD:B VSS:B
D1 VSS VDD diode_pd2nw_03v3 area='10u * 10u ' pj='2*10u + 2*10u ' m=4
.ends
