** sch_path: /foss/designs/libs/core_analog/pass1u05u/pass1u05u.sch
.subckt pass1u05u ind vss clkn ins clkp vdd
*.PININFO ind:B ins:B clkn:B clkp:B vdd:B vss:B
M1 ind clkp ins vdd pfet_03v3 L=0.5u W=3.0u nf=1 m=1
M2 ind clkn ins vss nfet_03v3 L=0.5u W=1.0u nf=1 m=1
.ends
