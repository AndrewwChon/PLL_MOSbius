** sch_path: /foss/designs/libs/qw_core_analog/SRegister_10/SRegister_10.sch
.include /foss/designs/switch_matrix_gf180mcu_9t5v0-main/gf180mcu_fd_sc_mcu9t5v0.spice
.subckt SRegister_10 VDDd VSSd phi1 phi2 en default[1] default[2] default[3] default[4] default[5] default[6] default[7]
+ default[8] default[9] default[10] d q out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8] out[9] out[10]
*.PININFO VDDd:B VSSd:B phi1:B phi2:B en:B default[1:10]:B d:B q:B out[1:10]:B
x11 net1 d phi1 phi2 VDDd VSSd out[1] en default[1] Register_unitcell
x1 net2 net1 phi1 phi2 VDDd VSSd out[2] en default[2] Register_unitcell
x2 net3 net2 phi1 phi2 VDDd VSSd out[3] en default[3] Register_unitcell
x3 net4 net3 phi1 phi2 VDDd VSSd out[4] en default[4] Register_unitcell
x4 net5 net4 phi1 phi2 VDDd VSSd out[5] en default[5] Register_unitcell
x5 net6 net5 phi1 phi2 VDDd VSSd out[6] en default[6] Register_unitcell
x6 net7 net6 phi1 phi2 VDDd VSSd out[7] en default[7] Register_unitcell
x7 net8 net7 phi1 phi2 VDDd VSSd out[8] en default[8] Register_unitcell
x8 net9 net8 phi1 phi2 VDDd VSSd out[9] en default[9] Register_unitcell
x9 q net9 phi1 phi2 VDDd VSSd out[10] en default[10] Register_unitcell
.ends

* expanding   symbol:  libs/qw_core_analog/Register_unitcell/Register_unitcell.sym # of pins=9
** sym_path: /foss/designs/libs/qw_core_analog/Register_unitcell/Register_unitcell.sym
** sch_path: /foss/designs/libs/qw_core_analog/Register_unitcell/Register_unitcell.sch
.subckt Register_unitcell q d phi1 phi2 VDDd VSSd out en default
*.PININFO phi1:B phi2:B d:B q:B en:B default:B out:B VDDd:B VSSd:B
x4 en enbar VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
* noconn VDDd
* noconn VSSd
x1 d q phi1 phi2 VDDd VSSd DFF_2phase_1
x2 q en or1 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1
x10 or2 or1 out VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1
x3 enbar default or2 VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1
.ends


* expanding   symbol:  libs/qw_core_analog/DFF_2phase_1/DFF_2phase_1.sym # of pins=6
** sym_path: /foss/designs/libs/qw_core_analog/DFF_2phase_1/DFF_2phase_1.sym
** sch_path: /foss/designs/libs/qw_core_analog/DFF_2phase_1/DFF_2phase_1.sch
.subckt DFF_2phase_1 D Q PHI_1 PHI_2 VDDd VSSd
*.PININFO D:I PHI_1:I PHI_2:I Q:O VDDd:B VSSd:B
* noconn VSSd
* noconn VDDd
xmain D PHI_1 out_m VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1
xsecondary out_m PHI_2 Q VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1
.ends

