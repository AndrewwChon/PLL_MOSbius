* NGSPICE file created from top_level_20250912_nosc.ext - technology: gf180mcuD

.subckt pfet a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$178 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$191 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$189 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$179 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$177 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$192 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0#
+ a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$190 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$180 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt asc_drive_buffer_up vss out in vdd
Xpfet_0 out out m1_778_712# vdd m1_778_712# out vdd vdd m1_778_712# out m1_778_712#
+ m1_778_712# out m1_778_712# vdd m1_778_712# vdd m1_778_712# pfet
Xpfet$178_0 vdd vdd m1_506_712# m1_n30_1318# pfet$178
Xnfet$191_0 m1_n566_1318# vss m1_n30_1318# vss nfet$191
Xnfet$189_0 out out vss m1_778_712# m1_778_712# out vss m1_778_712# m1_778_712# m1_778_712#
+ out m1_778_712# m1_778_712# out vss m1_778_712# vss vss nfet$189
Xpfet$179_0 vdd vdd m1_n30_1318# m1_n566_1318# pfet$179
Xpfet$177_0 m1_778_712# vdd vdd m1_778_712# m1_506_712# m1_506_712# m1_778_712# vdd
+ m1_506_712# m1_506_712# pfet$177
Xnfet$192_0 in vss m1_n566_1318# vss nfet$192
Xnfet_0 m1_778_712# vss m1_506_712# m1_506_712# m1_506_712# m1_778_712# m1_778_712#
+ vss m1_506_712# vss nfet
Xnfet$190_0 m1_n30_1318# vss m1_506_712# vss nfet$190
Xpfet$180_0 vdd vdd m1_n566_1318# in pfet$180
.ends

.subckt pfet$185 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$182 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$189 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$197 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$198 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$217 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$195 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$187 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$222 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$208 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$207 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$192 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$201 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$213 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$220 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$205 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$199 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$193 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$206 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$210 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$181 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$183 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$190 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$203 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$229 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$211 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$204 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$186 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$201 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$199 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$227 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$202 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$197 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$225 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$218 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$200 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$196 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$195 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$223 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$208 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$188 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$216 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$209 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$184 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$213 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$193 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$221 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$206 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$194 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$214 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$207 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$211 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$191 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$204 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$212 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$205 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$202 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$228 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$210 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$203 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$200 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$198 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$226 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$219 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$196 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$224 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$209 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$194 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$215 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$212 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt asc_dual_psd_def_20250809 vdd vss pd1 pd2 pd3 pd4 pd5 pd6 pd7 pd8 pd9 fout
+ sd1 sd2 sd3 sd4 sd5 sd6 sd7 sd8 sd9 fin define
Xpfet$185_17 vdd vdd m1_25739_21786# m1_25107_21786# pfet$185
Xpfet$182_108 vdd vdd m1_15454_18030# m1_15564_15778# pfet$182
Xpfet$189_6 vdd vdd m1_n290_24224# m1_n910_23922# pfet$189
Xnfet$197_5 m1_10458_17836# m1_11738_16080# m1_11271_18030# vss nfet$197
Xnfet$198_10 m1_21590_21786# vss m1_22222_21786# vss nfet$198
Xnfet$217_6 m1_27292_16202# m1_27292_16202# vss vss m1_26774_16398# vss nfet$217
Xnfet$195_2 m1_9288_21786# m1_9288_21786# m1_9645_21447# m1_9645_21447# m1_10509_21586#
+ vss nfet$195
Xpfet$187_3 vdd vdd m1_5901_19550# m1_649_17714# pfet$187
Xnfet$222_4 m1_n4978_24224# m1_n4978_24224# m1_n10452_25858# m1_n10452_25858# m1_n4880_24542#
+ vss nfet$222
Xnfet$208_2 m1_9645_21447# m1_9645_21447# vss vss m1_30492_21430# vss nfet$208
Xpfet$182_18 vdd m1_1119_17714# vdd m1_2194_16202# pfet$182
Xpfet$182_29 vdd vdd m1_1578_16080# m1_n7513_20152# pfet$182
Xpfet$207_4 vdd vdd m1_n5571_25662# m1_n10452_25858# pfet$207
Xpfet$192_1 vdd vdd m1_30256_19792# m1_21456_22513# pfet$192
Xnfet$201_9 m1_n10452_25858# vss m1_27031_17343# vss nfet$201
Xpfet$185_0 vdd vdd m1_n1133_21590# m1_n1263_21786# pfet$185
Xnfet$195_11 m1_19969_21590# m1_19969_21590# m1_21456_22513# m1_21456_22513# m1_20428_21586#
+ vss nfet$195
Xnfet$213_0 m1_7198_15778# m1_7198_15778# m1_7088_18030# m1_7088_18030# m1_7324_17358#
+ vss nfet$213
Xnfet$220_1 m1_n1927_20274# m1_n1927_20274# vss vss m1_n2445_20470# vss nfet$220
Xpfet$205_1 vdd m1_n8625_26174# vdd m1_n8848_25658# pfet$205
Xnfet$199_9 m1_25747_17714# vss m1_27003_19550# vss nfet$199
Xpfet$182_109 vdd vdd m1_10299_17343# m1_13198_17714# pfet$182
Xpfet$189_7 vdd vdd m1_32330_25662# m1_32193_25858# pfet$189
Xnfet$197_6 m1_6116_17343# vss m1_6275_17836# vss nfet$197
Xnfet$217_7 m1_26676_16080# m1_26676_16080# m1_26217_17714# m1_26217_17714# m1_26774_16398#
+ vss nfet$217
Xnfet$195_3 m1_9418_21590# m1_9418_21590# m1_9645_21447# m1_9645_21447# m1_9877_21586#
+ vss nfet$195
Xnfet$198_11 m1_18073_21786# vss m1_18705_21786# vss nfet$198
Xpfet$187_4 vdd vdd m1_12935_19550# m1_9015_17714# pfet$187
Xnfet$208_3 m1_7388_22513# m1_7388_22513# m1_30256_22102# m1_30256_22102# m1_30492_21430#
+ vss nfet$208
Xpfet$182_19 vdd m1_3015_15778# m1_2194_16202# m1_1933_17343# pfet$182
Xnfet$222_5 m1_n4362_24346# m1_n4362_24346# vss vss m1_n4880_24542# vss nfet$222
Xpfet$207_5 vdd vdd m1_n4847_25662# m1_n10452_25858# pfet$207
Xnfet$193_0 m1_4509_24346# m1_4509_24346# vss vss m1_3991_24542# vss nfet$193
Xpfet$192_2 vdd m1_30256_19792# vdd m1_24973_22513# pfet$192
Xpfet$185_1 vdd vdd m1_11671_21786# m1_11039_21786# pfet$185
Xnfet$195_12 m1_16322_21786# m1_16322_21786# m1_17939_22513# m1_17939_22513# m1_17543_21586#
+ vss nfet$195
Xnfet$213_1 m1_5761_16080# m1_5761_16080# vss vss m1_7324_17358# vss nfet$213
Xnfet$220_2 m1_n3206_20274# m1_n3206_20274# vss vss m1_n3724_20470# vss nfet$220
Xnfet$206_0 m1_11039_21786# m1_11039_21786# vss vss m1_9877_21586# vss nfet$206
Xpfet$205_2 vdd m1_n3651_26174# vdd m1_n4978_24224# pfet$205
Xpfet$210_0 vdd m1_n6380_21786# m1_n6380_21786# m1_n5019_19550# m1_n5227_20152# m1_n5227_20152#
+ pfet$210
Xnfet$197_7 m1_9485_17714# vss m1_10075_17518# vss nfet$197
Xpfet$189_8 vdd vdd m1_33174_24224# m1_32554_23922# pfet$189
Xpfet$181_110 vdd m1_11903_24542# vdd m1_12875_24346# pfet$181
Xnfet$198_12 m1_14556_21786# vss m1_15188_21786# vss nfet$198
Xpfet$187_5 vdd vdd m1_8137_20152# m1_965_15478# pfet$187
Xnfet$195_4 m1_5901_21590# m1_5901_21590# m1_7388_22513# m1_7388_22513# m1_6360_21586#
+ vss nfet$195
Xnfet$222_6 m1_n4978_24224# m1_n4978_24224# vss vss m1_n3415_25502# vss nfet$222
Xnfet$193_1 m1_3893_24224# m1_3893_24224# m1_3537_24542# m1_3537_24542# m1_3991_24542#
+ vss nfet$193
Xpfet$192_3 vdd vdd m1_34843_21786# m1_34093_19792# pfet$192
Xpfet$207_6 vdd vdd m1_n4623_25487# fin pfet$207
Xpfet$185_2 vdd vdd m1_12935_21590# m1_12805_21786# pfet$185
Xnfet$195_13 m1_16452_21590# m1_16452_21590# m1_17939_22513# m1_17939_22513# m1_16911_21586#
+ vss nfet$195
Xnfet$213_2 m1_9944_16080# m1_9944_16080# vss vss m1_11507_17358# vss nfet$213
Xnfet$220_3 m1_n6973_21481# m1_n6973_21481# m1_n6839_20152# m1_n6839_20152# m1_n6282_20470#
+ vss nfet$220
Xpfet$205_3 vdd vdd m1_n3651_26174# m1_n3541_23922# pfet$205
Xnfet$206_1 m1_11671_21786# m1_11671_21786# vss vss m1_10509_21586# vss nfet$206
Xpfet$183_30 vdd vdd vdd m1_17539_22402# m1_16322_21786# m1_16322_21786# pfet$183
Xpfet$190_0 vdd vdd m1_n646_24542# m1_n290_24224# pfet$190
Xpfet$210_1 vdd vdd vdd m1_n5019_22344# m1_n4485_21904# m1_n4485_21904# pfet$210
Xpfet$203_0 vdd m1_n10309_25662# m1_n10572_23922# m1_n10796_25662# pfet$203
Xnfet$201_10 m1_26217_17714# vss m1_29087_15778# vss nfet$201
Xnfet$197_8 m1_7555_16080# vss m1_7198_15778# vss nfet$197
Xpfet$189_9 vdd vdd m1_28624_21786# m1_32675_25947# pfet$189
Xpfet$181_100 vdd vdd m1_29607_24346# m1_n7513_20152# pfet$181
Xnfet$198_13 m1_16322_21786# vss m1_16452_21590# vss nfet$198
Xnfet$229_0 m1_n6839_20152# vss m1_n8145_21908# vss nfet$229
Xnfet$195_5 m1_2254_21786# m1_2254_21786# m1_3871_22513# m1_3871_22513# m1_3475_21586#
+ vss nfet$195
Xpfet$187_6 vdd vdd m1_9418_19550# m1_4832_17714# pfet$187
Xnfet$193_2 m1_4997_25658# m1_4997_25658# vss vss m1_5456_25502# vss nfet$193
Xnfet$222_7 m1_n3541_23922# m1_n3541_23922# m1_n3651_26174# m1_n3651_26174# m1_n3415_25502#
+ vss nfet$222
Xpfet$192_4 vdd m1_34093_19792# vdd m1_32818_20470# pfet$192
Xpfet$207_7 vdd vdd m1_n3541_23922# m1_n3184_24224# pfet$207
Xpfet$185_3 vdd vdd m1_9418_21590# m1_9288_21786# pfet$185
Xnfet$195_14 m1_12805_21786# m1_12805_21786# m1_14422_22513# m1_14422_22513# m1_14026_21586#
+ vss nfet$195
Xnfet$213_3 m1_11381_15778# m1_11381_15778# m1_11271_18030# m1_11271_18030# m1_11507_17358#
+ vss nfet$213
Xnfet$220_4 m1_2590_19404# m1_2590_19404# vss vss m1_n2445_21430# vss nfet$220
Xnfet$206_2 m1_8154_21786# m1_8154_21786# vss vss m1_6992_21586# vss nfet$206
Xpfet$183_31 vdd vdd vdd m1_27462_22102# m1_27003_21590# m1_27003_21590# pfet$183
Xpfet$183_20 vdd vdd vdd m1_20428_22102# m1_19969_21590# m1_19969_21590# pfet$183
Xpfet$190_1 vdd m1_n789_25858# vdd m1_814_25658# pfet$190
Xpfet$183_0 vdd vdd vdd m1_n674_22102# m1_n1133_21590# m1_n1133_21590# pfet$183
Xpfet$205_4 vdd m1_n10452_25858# vdd m1_n4362_24346# pfet$205
Xnfet$211_0 m1_34093_22102# vss fout vss nfet$211
Xpfet$210_2 vdd m1_n5764_21786# m1_n5764_21786# m1_n5019_22344# m1_n5227_21418# m1_n5227_21418#
+ pfet$210
Xpfet$203_1 vdd m1_n9952_24224# m1_n8848_25658# m1_n10933_25858# pfet$203
Xnfet$201_11 m1_27031_17343# vss m1_27190_17836# vss nfet$201
Xnfet$197_9 sd5 vss m1_9331_15478# vss nfet$197
Xpfet$181_101 vdd vdd m1_28010_25858# m1_21590_21786# pfet$181
Xnfet$198_14 m1_19839_21786# vss m1_19969_21590# vss nfet$198
Xnfet$195_6 m1_2384_21590# m1_2384_21590# m1_3871_22513# m1_3871_22513# m1_2843_21586#
+ vss nfet$195
Xpfet$187_7 vdd vdd m1_11654_20152# m1_5148_15478# pfet$187
Xpfet$192_5 vdd vdd m1_34093_19792# m1_32818_21586# pfet$192
Xnfet$193_3 m1_4509_24346# m1_4509_24346# m1_3394_25858# m1_3394_25858# m1_5456_25502#
+ vss nfet$193
Xpfet$207_8 vdd vdd m1_n2567_23922# m1_n7320_25516# pfet$207
Xpfet$185_4 vdd vdd m1_8154_21786# m1_7522_21786# pfet$185
Xnfet$195_15 m1_26873_21786# m1_26873_21786# m1_28490_22513# m1_28490_22513# m1_28094_21586#
+ vss nfet$195
Xnfet$213_4 m1_10560_16202# m1_10560_16202# vss vss m1_10042_16398# vss nfet$213
Xnfet$220_5 m1_6107_19404# m1_6107_19404# m1_n5227_21418# m1_n5227_21418# m1_n2445_21430#
+ vss nfet$220
Xnfet$206_3 m1_7522_21786# m1_7522_21786# vss vss m1_6360_21586# vss nfet$206
Xpfet$183_32 vdd m1_28490_22513# m1_28490_22513# m1_28090_22402# m1_28624_21786# m1_28624_21786#
+ pfet$183
Xpfet$183_21 vdd vdd vdd m1_21056_22402# m1_19839_21786# m1_19839_21786# pfet$183
Xpfet$190_2 vdd vdd m1_n789_25858# m1_326_24346# pfet$190
Xpfet$205_5 vdd vdd m1_n10308_24542# m1_n9952_24224# pfet$205
Xpfet$183_1 vdd m1_7388_22513# m1_7388_22513# m1_6988_22402# m1_7522_21786# m1_7522_21786#
+ pfet$183
Xpfet$183_10 vdd m1_3871_22513# m1_3871_22513# m1_2843_22102# m1_4637_21786# m1_4637_21786#
+ pfet$183
Xnfet$204_0 pd1 vss m1_n1263_21786# vss nfet$204
Xpfet$203_2 vdd m1_n4362_24346# m1_n4847_25662# m1_n4464_25980# pfet$203
Xnfet$201_12 m1_28470_16080# vss m1_28113_15778# vss nfet$201
Xpfet$181_102 vdd m1_28371_23922# m1_28635_24542# m1_28010_25858# pfet$181
Xnfet$198_15 m1_28624_21786# vss m1_29256_21786# vss nfet$198
Xnfet$195_7 m1_5771_21786# m1_5771_21786# m1_7388_22513# m1_7388_22513# m1_6992_21586#
+ vss nfet$195
Xpfet$187_8 vdd vdd m1_n1133_19550# m1_n7383_17599# pfet$187
Xpfet$186_10 vdd vdd m1_27031_17343# m1_n10452_25858# pfet$186
Xnfet$193_4 m1_12259_24224# m1_12259_24224# m1_11903_24542# m1_11903_24542# m1_12357_24542#
+ vss nfet$193
Xpfet$207_9 vdd vdd m1_n4464_25980# m1_n4623_25487# pfet$207
Xpfet$192_6 vdd vdd m1_31535_19792# m1_14422_22513# pfet$192
Xpfet$185_5 vdd vdd m1_1120_21786# m1_488_21786# pfet$185
Xnfet$195_16 m1_27003_21590# m1_27003_21590# m1_28490_22513# m1_28490_22513# m1_27462_21586#
+ vss nfet$195
Xnfet$213_5 m1_9944_16080# m1_9944_16080# m1_9485_17714# m1_9485_17714# m1_10042_16398#
+ vss nfet$213
Xnfet$220_6 m1_n5764_21786# m1_n5764_21786# vss vss m1_n6282_21430# vss nfet$220
Xnfet$206_4 m1_1120_21786# m1_1120_21786# vss vss m1_n42_21586# vss nfet$206
Xpfet$190_3 vdd m1_n646_24542# vdd m1_326_24346# pfet$190
Xpfet$205_6 vdd m1_n10308_24542# vdd m1_n9336_24346# pfet$205
Xpfet$183_2 vdd m1_7388_22513# m1_7388_22513# m1_6360_22102# m1_8154_21786# m1_8154_21786#
+ pfet$183
Xpfet$183_33 vdd m1_28490_22513# m1_28490_22513# m1_27462_22102# m1_29256_21786# m1_29256_21786#
+ pfet$183
Xpfet$183_22 vdd m1_21456_22513# m1_21456_22513# m1_20428_22102# m1_22222_21786# m1_22222_21786#
+ pfet$183
Xpfet$183_11 vdd vdd vdd m1_2843_22102# m1_2384_21590# m1_2384_21590# pfet$183
Xnfet$204_1 pd2 vss m1_2254_21786# vss nfet$204
Xpfet$203_3 vdd m1_n3184_24224# m1_n3651_26174# m1_n4623_25487# pfet$203
Xnfet$201_13 m1_26217_17714# vss m1_25747_17714# vss nfet$201
Xpfet$189_10 vdd vdd m1_35071_24542# m1_32675_25947# pfet$189
Xpfet$201_0 vdd vdd m1_n7513_20152# m1_35837_22102# pfet$201
Xpfet$181_103 vdd vdd m1_28635_24542# m1_28991_24224# pfet$181
Xnfet$195_8 m1_23486_21590# m1_23486_21590# m1_24973_22513# m1_24973_22513# m1_23945_21586#
+ vss nfet$195
Xnfet$198_16 m1_26873_21786# vss m1_27003_21590# vss nfet$198
Xpfet$187_9 vdd vdd m1_27003_19550# m1_25747_17714# pfet$187
Xpfet$186_11 vdd vdd m1_26807_17518# m1_26217_17714# pfet$186
Xpfet$199_0 vdd vdd m1_n7247_17714# m1_n6788_16080# pfet$199
Xnfet$193_5 m1_8692_24346# m1_8692_24346# vss vss m1_8174_24542# vss nfet$193
Xpfet$192_7 vdd vdd m1_31535_22102# m1_354_22513# pfet$192
Xnfet$227_0 m1_n927_19404# m1_n927_19404# vss vss m1_n6282_20470# vss nfet$227
Xpfet$185_6 vdd vdd m1_5901_21590# m1_5771_21786# pfet$185
Xnfet$195_17 m1_12935_21590# m1_12935_21590# m1_14422_22513# m1_14422_22513# m1_13394_21586#
+ vss nfet$195
Xnfet$213_6 m1_1578_16080# m1_1578_16080# vss vss m1_3141_17358# vss nfet$213
Xnfet$220_7 m1_n3822_21786# m1_n3822_21786# m1_n4485_21904# m1_n4485_21904# m1_n3724_21430#
+ vss nfet$220
Xnfet$206_5 m1_4005_21786# m1_4005_21786# vss vss m1_2843_21586# vss nfet$206
Xpfet$190_4 vdd vdd m1_32675_25947# m1_33790_24346# pfet$190
Xpfet$205_7 vdd vdd m1_n10452_25858# m1_n4978_24224# pfet$205
Xpfet$183_3 vdd m1_9645_21447# m1_9645_21447# m1_10505_22402# m1_11039_21786# m1_11039_21786#
+ pfet$183
Xpfet$183_34 vdd vdd vdd m1_28090_22402# m1_26873_21786# m1_26873_21786# pfet$183
Xpfet$183_23 vdd vdd vdd m1_23945_22102# m1_23486_21590# m1_23486_21590# pfet$183
Xpfet$183_12 vdd vdd vdd m1_3471_22402# m1_2254_21786# m1_2254_21786# pfet$183
Xnfet$204_2 pd9 vss m1_26873_21786# vss nfet$204
Xpfet$203_4 vdd m1_n2567_23922# m1_n3184_24224# m1_n4464_25980# pfet$203
Xpfet$181_0 vdd vdd m1_3049_25662# m1_2912_25858# pfet$181
Xpfet$189_11 vdd vdd m1_32817_25662# m1_32675_25947# pfet$189
Xpfet$181_104 vdd m1_25912_25658# m1_26705_24542# m1_23964_25662# pfet$181
Xnfet$198_17 m1_25107_21786# vss m1_25739_21786# vss nfet$198
Xnfet$195_9 m1_23356_21786# m1_23356_21786# m1_24973_22513# m1_24973_22513# m1_24577_21586#
+ vss nfet$195
Xpfet$186_12 vdd vdd m1_26676_16080# m1_n7513_20152# pfet$186
Xpfet$199_1 vdd m1_n7247_17714# vdd m1_n6172_16202# pfet$199
Xnfet$193_6 m1_8076_24224# m1_8076_24224# m1_7720_24542# m1_7720_24542# m1_8174_24542#
+ vss nfet$193
Xnfet$227_1 m1_n2543_20130# m1_n2543_20130# m1_n5227_20152# m1_n5227_20152# m1_n2445_20470#
+ vss nfet$227
Xpfet$185_7 vdd vdd m1_4637_21786# m1_4005_21786# pfet$185
Xnfet$213_7 m1_5761_16080# m1_5761_16080# m1_5302_17714# m1_5302_17714# m1_5859_16398#
+ vss nfet$213
Xnfet$220_8 m1_9624_19404# m1_9624_19404# vss vss m1_n3724_21430# vss nfet$220
Xnfet$206_6 m1_4637_21786# m1_4637_21786# vss vss m1_3475_21586# vss nfet$206
Xpfet$183_35 vdd vdd vdd m1_13394_22102# m1_12935_21590# m1_12935_21590# pfet$183
Xpfet$190_5 vdd m1_32675_25947# vdd m1_34278_25658# pfet$190
Xpfet$183_24 vdd m1_17939_22513# m1_17939_22513# m1_16911_22102# m1_18705_21786# m1_18705_21786#
+ pfet$183
Xpfet$183_13 vdd vdd vdd m1_6988_22402# m1_5771_21786# m1_5771_21786# pfet$183
Xpfet$183_4 vdd vdd vdd m1_9877_22102# m1_9418_21590# m1_9418_21590# pfet$183
Xpfet$181_1 vdd m1_3536_25662# m1_3273_23922# m1_3049_25662# pfet$181
Xpfet$203_5 vdd m1_n10572_23922# m1_n10308_24542# m1_n10933_25858# pfet$203
Xnfet$202_0 m1_n10452_25858# vss m1_n1271_25858# vss nfet$202
Xpfet$189_12 vdd vdd m1_32193_25858# m1_25107_21786# pfet$189
Xpfet$181_105 vdd vdd m1_30888_24542# m1_28492_25858# pfet$181
Xpfet$181_90 vdd vdd m1_24309_25858# m1_25424_24346# pfet$181
Xpfet$199_2 vdd vdd m1_n5461_18030# m1_n5351_15778# pfet$199
Xpfet$186_13 vdd vdd m1_25747_17714# m1_26217_17714# pfet$186
Xnfet$193_7 m1_9180_25658# m1_9180_25658# vss vss m1_9639_25502# vss nfet$193
Xpfet$185_8 vdd vdd m1_2384_21590# m1_2254_21786# pfet$185
Xnfet$206_7 m1_488_21786# m1_488_21786# vss vss m1_n674_21586# vss nfet$206
Xnfet$213_8 m1_3015_15778# m1_3015_15778# m1_2905_18030# m1_2905_18030# m1_3141_17358#
+ vss nfet$213
Xnfet$220_9 m1_n6380_21786# m1_n6380_21786# m1_n6839_21786# m1_n6839_21786# m1_n6282_21430#
+ vss nfet$220
Xpfet$190_6 vdd vdd m1_32818_24542# m1_33174_24224# pfet$190
Xpfet$183_25 vdd m1_17939_22513# m1_17939_22513# m1_17539_22402# m1_18073_21786# m1_18073_21786#
+ pfet$183
Xpfet$183_14 vdd vdd vdd m1_n46_22402# m1_n1263_21786# m1_n1263_21786# pfet$183
Xpfet$183_5 vdd m1_9645_21447# m1_9645_21447# m1_9877_22102# m1_11671_21786# m1_11671_21786#
+ pfet$183
Xpfet$181_2 vdd vdd m1_3394_25858# m1_4509_24346# pfet$181
Xpfet$203_6 vdd m1_n8848_25658# m1_n8055_24542# m1_n10796_25662# pfet$203
Xnfet$202_1 m1_n789_25858# vss m1_n647_25662# vss nfet$202
Xpfet$189_13 vdd vdd m1_33790_24346# m1_n7513_20152# pfet$189
Xpfet$181_106 vdd vdd m1_25107_21786# m1_28492_25858# pfet$181
Xpfet$181_91 vdd vdd m1_23356_21786# pd8 pfet$181
Xpfet$181_80 vdd vdd m1_17058_24346# m1_n7513_20152# pfet$181
Xpfet$199_3 vdd m1_n5461_18030# vdd m1_n6788_16080# pfet$199
Xpfet$185_9 vdd vdd m1_22222_21786# m1_21590_21786# pfet$185
Xnfet$193_8 m1_8692_24346# m1_8692_24346# m1_7577_25858# m1_7577_25858# m1_9639_25502#
+ vss nfet$193
Xpfet$197_0 vdd vdd fout m1_34093_22102# pfet$197
Xnfet$206_8 m1_25739_21786# m1_25739_21786# vss vss m1_24577_21586# vss nfet$206
Xnfet$213_9 m1_2194_16202# m1_2194_16202# vss vss m1_1676_16398# vss nfet$213
Xpfet$190_7 vdd m1_32818_24542# vdd m1_33790_24346# pfet$190
Xpfet$183_26 vdd vdd vdd m1_16911_22102# m1_16452_21590# m1_16452_21590# pfet$183
Xpfet$183_15 vdd m1_354_22513# m1_354_22513# m1_n46_22402# m1_488_21786# m1_488_21786#
+ pfet$183
Xnfet$225_0 m1_n8283_20611# vss m1_n8283_19850# vss nfet$225
Xpfet$183_6 vdd vdd vdd m1_10505_22402# m1_9288_21786# m1_9288_21786# pfet$183
Xpfet$203_7 vdd m1_n3541_23922# m1_n4362_24346# m1_n4623_25487# pfet$203
Xpfet$181_3 vdd m1_3394_25858# vdd m1_4997_25658# pfet$181
Xnfet$202_2 m1_n1271_25858# vss m1_n1134_25662# vss nfet$202
Xpfet$181_107 vdd m1_24309_25858# vdd m1_25912_25658# pfet$181
Xnfet$193_20 m1_21241_24346# m1_21241_24346# m1_20126_25858# m1_20126_25858# m1_22188_25502#
+ vss nfet$193
Xpfet$181_92 vdd vdd m1_28492_25858# m1_29607_24346# pfet$181
Xpfet$181_81 vdd vdd m1_18339_24542# m1_15943_25858# pfet$181
Xpfet$181_70 vdd vdd m1_14156_24542# m1_11760_25858# pfet$181
Xpfet$199_4 vdd vdd m1_26217_17714# m1_26676_16080# pfet$199
Xnfet$193_9 m1_17058_24346# m1_17058_24346# vss vss m1_16540_24542# vss nfet$193
Xnfet$206_9 m1_25107_21786# m1_25107_21786# vss vss m1_23945_21586# vss nfet$206
Xnfet$225_1 m1_n7513_20152# m1_n8283_19850# vss vss nfet$225
Xnfet$218_0 m1_n10452_25858# m1_n10452_25858# m1_n7186_25858# m1_n7186_25858# m1_n6629_25502#
+ vss nfet$218
Xpfet$183_7 vdd m1_354_22513# m1_354_22513# m1_n674_22102# m1_1120_21786# m1_1120_21786#
+ pfet$183
Xpfet$183_27 vdd m1_14422_22513# m1_14422_22513# m1_14022_22402# m1_14556_21786# m1_14556_21786#
+ pfet$183
Xpfet$183_16 vdd m1_24973_22513# m1_24973_22513# m1_23945_22102# m1_25739_21786# m1_25739_21786#
+ pfet$183
Xpfet$181_4 vdd vdd m1_3893_24224# m1_3273_23922# pfet$181
Xnfet$202_3 m1_n7513_20152# vss m1_326_24346# vss nfet$202
Xpfet$181_108 vdd vdd m1_25424_24346# m1_n7513_20152# pfet$181
Xnfet$193_21 m1_28991_24224# m1_28991_24224# m1_28635_24542# m1_28635_24542# m1_29089_24542#
+ vss nfet$193
Xnfet$193_10 m1_17546_25658# m1_17546_25658# vss vss m1_18005_25502# vss nfet$193
Xnfet$200_0 sd9 vss m1_n7401_15478# vss nfet$200
Xpfet$181_93 vdd m1_28991_24224# m1_30095_25658# m1_28010_25858# pfet$181
Xpfet$181_82 vdd vdd m1_21241_24346# m1_n7513_20152# pfet$181
Xpfet$181_71 vdd vdd m1_11039_21786# m1_11760_25858# pfet$181
Xpfet$181_60 vdd vdd m1_20126_25858# m1_21241_24346# pfet$181
Xpfet$199_5 vdd m1_26217_17714# vdd m1_27292_16202# pfet$199
Xnfet$198_0 m1_n1263_21786# vss m1_n1133_21590# vss nfet$198
Xnfet$225_2 m1_n8145_21908# vss m1_n8283_20611# vss nfet$225
Xnfet$218_1 m1_n6111_25858# m1_n6111_25858# vss vss m1_n6629_25502# vss nfet$218
Xpfet$183_8 vdd vdd vdd m1_6360_22102# m1_5901_21590# m1_5901_21590# pfet$183
Xpfet$183_28 vdd m1_14422_22513# m1_14422_22513# m1_13394_22102# m1_15188_21786# m1_15188_21786#
+ pfet$183
Xpfet$183_17 vdd m1_21456_22513# m1_21456_22513# m1_21056_22402# m1_21590_21786# m1_21590_21786#
+ pfet$183
Xnfet$196_10 m1_9015_17714# m1_9015_17714# vss vss m1_14005_20470# vss nfet$196
Xpfet$181_5 vdd m1_3893_24224# m1_4997_25658# m1_2912_25858# pfet$181
Xnfet$202_4 m1_n789_25858# vss m1_1607_24542# vss nfet$202
Xpfet$181_109 vdd m1_12259_24224# m1_13363_25658# m1_11278_25858# pfet$181
Xnfet$193_22 m1_29607_24346# m1_29607_24346# vss vss m1_29089_24542# vss nfet$193
Xnfet$193_11 m1_16442_24224# m1_16442_24224# m1_16086_24542# m1_16086_24542# m1_16540_24542#
+ vss nfet$193
Xnfet$200_1 sd2 vss m1_21880_15478# vss nfet$200
Xpfet$181_94 vdd m1_28492_25858# vdd m1_30095_25658# pfet$181
Xpfet$181_83 vdd m1_21729_25658# m1_22522_24542# m1_19781_25662# pfet$181
Xpfet$181_72 vdd m1_13363_25658# m1_14156_24542# m1_11415_25662# pfet$181
Xpfet$181_61 vdd m1_24452_24542# vdd m1_25424_24346# pfet$181
Xpfet$181_50 vdd vdd m1_20268_25662# m1_20126_25858# pfet$181
Xpfet$199_6 vdd vdd m1_28003_18030# m1_28113_15778# pfet$199
Xnfet$199_10 m1_26063_15478# vss m1_29239_20152# vss nfet$199
Xnfet$198_1 m1_11039_21786# vss m1_11671_21786# vss nfet$198
Xnfet$225_3 m1_n8283_19850# m1_n8283_20611# vss vss nfet$225
Xpfet$195_0 vdd m1_34093_22102# vdd m1_28490_22513# pfet$195
Xpfet$183_29 vdd vdd vdd m1_14022_22402# m1_12805_21786# m1_12805_21786# pfet$183
Xpfet$183_18 vdd vdd vdd m1_24573_22402# m1_23356_21786# m1_23356_21786# pfet$183
Xpfet$183_9 vdd m1_3871_22513# m1_3871_22513# m1_3471_22402# m1_4005_21786# m1_4005_21786#
+ pfet$183
Xnfet$196_11 m1_13198_17714# m1_13198_17714# vss vss m1_17522_20470# vss nfet$196
Xpfet$181_6 vdd vdd m1_3536_25662# m1_3394_25858# pfet$181
Xnfet$223_0 m1_n10933_25858# m1_n8848_25658# m1_n8055_24542# vss nfet$223
Xpfet$208_0 vdd vdd m1_n7186_25858# m1_n10452_25858# pfet$208
Xnfet$202_5 m1_n789_25858# vss m1_488_21786# vss nfet$202
Xnfet$200_2 sd1 vss m1_26063_15478# vss nfet$200
Xnfet$193_23 m1_25424_24346# m1_25424_24346# m1_24309_25858# m1_24309_25858# m1_26371_25502#
+ vss nfet$193
Xnfet$193_12 m1_17058_24346# m1_17058_24346# m1_15943_25858# m1_15943_25858# m1_18005_25502#
+ vss nfet$193
Xpfet$181_95 vdd vdd m1_28991_24224# m1_28371_23922# pfet$181
Xpfet$181_84 vdd vdd m1_23827_25858# m1_18073_21786# pfet$181
Xpfet$181_73 vdd m1_16086_24542# vdd m1_17058_24346# pfet$181
Xpfet$181_62 vdd vdd m1_24452_24542# m1_24808_24224# pfet$181
Xpfet$181_51 vdd vdd m1_20625_24224# m1_20005_23922# pfet$181
Xpfet$181_40 vdd vdd m1_11760_25858# m1_12875_24346# pfet$181
Xpfet$199_7 vdd m1_28003_18030# vdd m1_26676_16080# pfet$199
Xnfet$199_11 m1_9331_15478# vss m1_15171_20152# vss nfet$199
Xnfet$198_2 m1_12805_21786# vss m1_12935_21590# vss nfet$198
Xpfet$183_19 vdd m1_24973_22513# m1_24973_22513# m1_24573_22402# m1_25107_21786# m1_25107_21786#
+ pfet$183
Xpfet$195_1 vdd vdd m1_34093_22102# m1_34843_21786# pfet$195
Xpfet$188_0 vdd vdd m1_n7401_15478# sd9 pfet$188
Xnfet$196_12 m1_16452_19550# m1_16452_19550# vss vss m1_16890_20470# vss nfet$196
Xpfet$181_7 vdd vdd m1_7232_25662# m1_7095_25858# pfet$181
Xnfet$216_0 m1_n6274_17836# m1_n4994_16080# m1_n5461_18030# vss nfet$216
Xnfet$223_1 m1_n10796_25662# m1_n10572_23922# m1_n10308_24542# vss nfet$223
Xpfet$208_1 vdd m1_n7186_25858# vdd m1_n6111_25858# pfet$208
Xnfet$202_6 m1_n910_23922# vss m1_n290_24224# vss nfet$202
Xnfet$193_24 m1_30095_25658# m1_30095_25658# vss vss m1_30554_25502# vss nfet$193
Xnfet$193_13 m1_13363_25658# m1_13363_25658# vss vss m1_13822_25502# vss nfet$193
Xpfet$181_96 vdd m1_28635_24542# vdd m1_29607_24346# pfet$181
Xpfet$181_85 vdd m1_24188_23922# m1_24452_24542# m1_23827_25858# pfet$181
Xpfet$181_74 vdd vdd m1_14556_21786# m1_15943_25858# pfet$181
Xpfet$181_63 vdd vdd m1_19781_25662# m1_19644_25858# pfet$181
Xpfet$181_52 vdd m1_20268_25662# m1_20005_23922# m1_19781_25662# pfet$181
Xpfet$181_41 vdd vdd m1_9288_21786# pd4 pfet$181
Xpfet$181_30 vdd vdd m1_2912_25858# m1_488_21786# pfet$181
Xnfet$199_12 m1_13514_15478# vss m1_18688_20152# vss nfet$199
Xnfet$198_3 m1_9288_21786# vss m1_9418_21590# vss nfet$198
Xnfet$196_0 m1_n3534_17714# m1_n3534_17714# vss vss m1_3454_20470# vss nfet$196
Xpfet$195_2 vdd vdd m1_30256_22102# m1_7388_22513# pfet$195
Xpfet$188_1 vdd vdd m1_21880_15478# sd2 pfet$188
Xnfet$196_13 m1_19969_19550# m1_19969_19550# vss vss m1_20407_20470# vss nfet$196
Xnfet$223_2 m1_n10933_25858# m1_n10309_25662# m1_n10572_23922# vss nfet$223
Xnfet$209_0 m1_31535_22102# m1_32818_21586# vss vss nfet$209
Xpfet$181_8 vdd vdd m1_8076_24224# m1_7456_23922# pfet$181
Xnfet$216_1 m1_n6433_17343# m1_n4377_15778# m1_n4994_16080# vss nfet$216
Xnfet$202_7 m1_25107_21786# vss m1_32193_25858# vss nfet$202
Xpfet$184_30 vdd vdd vdd m1_24560_19550# m1_21880_15478# m1_21880_15478# pfet$184
Xpfet$213_0 vdd vdd m1_n8145_21908# m1_n6839_20152# pfet$213
Xnfet$193_25 m1_29607_24346# m1_29607_24346# m1_28492_25858# m1_28492_25858# m1_30554_25502#
+ vss nfet$193
Xnfet$193_14 m1_12875_24346# m1_12875_24346# m1_11760_25858# m1_11760_25858# m1_13822_25502#
+ vss nfet$193
Xnfet$202_10 m1_32675_25947# vss m1_35071_24542# vss nfet$202
Xpfet$181_97 vdd vdd m1_21590_21786# m1_24309_25858# pfet$181
Xpfet$181_86 vdd m1_28634_25662# m1_28371_23922# m1_28147_25662# pfet$181
Xpfet$181_75 vdd vdd m1_19644_25858# m1_14556_21786# pfet$181
Xpfet$181_64 vdd vdd m1_22522_24542# m1_20126_25858# pfet$181
Xpfet$181_53 vdd m1_20625_24224# m1_21729_25658# m1_19644_25858# pfet$181
Xpfet$181_42 vdd m1_11760_25858# vdd m1_13363_25658# pfet$181
Xpfet$181_31 vdd m1_3273_23922# m1_3537_24542# m1_2912_25858# pfet$181
Xpfet$181_20 vdd vdd m1_4509_24346# m1_n7513_20152# pfet$181
Xnfet$213_20 m1_22493_16080# m1_22493_16080# m1_22034_17714# m1_22034_17714# m1_22591_16398#
+ vss nfet$213
Xnfet$199_13 m1_13198_17714# vss m1_16452_19550# vss nfet$199
Xnfet$198_4 m1_7522_21786# vss m1_8154_21786# vss nfet$198
Xnfet$196_1 m1_2384_19550# m1_2384_19550# vss vss m1_2822_20470# vss nfet$196
Xpfet$188_2 vdd vdd m1_26063_15478# sd1 pfet$188
Xpfet$195_3 vdd m1_31535_22102# vdd m1_3871_22513# pfet$195
Xnfet$196_14 m1_17381_17714# m1_17381_17714# vss vss m1_21039_20470# vss nfet$196
Xpfet$181_9 vdd m1_7719_25662# m1_7456_23922# m1_7232_25662# pfet$181
Xnfet$216_2 m1_n6274_17836# m1_n5351_15778# m1_n6172_16202# vss nfet$216
Xnfet$223_3 m1_n10796_25662# m1_n9952_24224# m1_n8848_25658# vss nfet$223
Xpfet$184_31 vdd m1_n2543_20130# m1_n2543_20130# m1_20407_19850# m1_19969_19550# m1_19969_19550#
+ pfet$184
Xpfet$184_20 vdd m1_n3822_21786# m1_n3822_21786# m1_14009_19550# m1_9015_17714# m1_9015_17714#
+ pfet$184
Xpfet$193_0 vdd m1_n647_25662# m1_n910_23922# m1_n1134_25662# pfet$193
Xnfet$202_8 m1_32193_25858# vss m1_32330_25662# vss nfet$202
Xnfet$221_0 m1_n8625_26174# vss m1_n8055_24542# vss nfet$221
Xpfet$206_0 vdd vdd m1_n4485_20152# m1_n3822_20130# pfet$206
Xnfet$193_26 m1_25912_25658# m1_25912_25658# vss vss m1_26371_25502# vss nfet$193
Xnfet$193_15 m1_25424_24346# m1_25424_24346# vss vss m1_24906_24542# vss nfet$193
Xnfet$202_11 m1_32554_23922# vss m1_33174_24224# vss nfet$202
Xpfet$181_98 vdd m1_30095_25658# m1_30888_24542# m1_28147_25662# pfet$181
Xpfet$181_87 vdd vdd m1_28147_25662# m1_28010_25858# pfet$181
Xpfet$181_76 vdd m1_20005_23922# m1_20269_24542# m1_19644_25858# pfet$181
Xpfet$181_65 vdd vdd m1_18073_21786# m1_20126_25858# pfet$181
Xpfet$181_54 vdd vdd m1_24808_24224# m1_24188_23922# pfet$181
Xpfet$181_43 vdd vdd m1_12805_21786# pd5 pfet$181
Xpfet$181_32 vdd vdd m1_7720_24542# m1_8076_24224# pfet$181
Xpfet$181_21 vdd m1_7456_23922# m1_7720_24542# m1_7095_25858# pfet$181
Xpfet$181_10 vdd m1_8076_24224# m1_9180_25658# m1_7095_25858# pfet$181
Xnfet$194_80 m1_28147_25662# m1_28991_24224# m1_30095_25658# vss nfet$194
Xnfet$213_21 m1_14127_16080# m1_14127_16080# vss vss m1_15690_17358# vss nfet$213
Xnfet$213_10 m1_1578_16080# m1_1578_16080# m1_1119_17714# m1_1119_17714# m1_1676_16398#
+ vss nfet$213
Xnfet$199_14 m1_21564_17714# vss m1_23486_19550# vss nfet$199
Xnfet$198_5 m1_488_21786# vss m1_1120_21786# vss nfet$198
Xpfet$195_4 vdd m1_30256_22102# vdd m1_9645_21447# pfet$195
Xnfet$196_2 m1_5901_19550# m1_5901_19550# vss vss m1_6339_20470# vss nfet$196
Xnfet$196_15 m1_21564_17714# m1_21564_17714# vss vss m1_24556_20470# vss nfet$196
Xnfet$216_3 m1_n6433_17343# m1_n6172_16202# m1_n6657_17518# vss nfet$216
Xnfet$223_4 m1_n4623_25487# m1_n2567_23922# m1_n3184_24224# vss nfet$223
Xpfet$184_32 vdd m1_n2543_20130# m1_n2543_20130# m1_21043_19550# m1_17381_17714# m1_17381_17714#
+ pfet$184
Xpfet$184_21 vdd vdd vdd m1_13373_19850# m1_15171_20152# m1_15171_20152# pfet$184
Xpfet$184_10 vdd vdd vdd m1_9856_19850# m1_11654_20152# m1_11654_20152# pfet$184
Xpfet$186_0 vdd vdd m1_n6274_17836# m1_n6433_17343# pfet$186
Xnfet$221_10 vss vss m1_n4978_24224# vss nfet$221
Xpfet$193_1 vdd m1_n910_23922# m1_n646_24542# m1_n1271_25858# pfet$193
Xnfet$202_9 m1_n7513_20152# vss m1_33790_24346# vss nfet$202
Xnfet$197_80 m1_18824_17836# m1_19747_15778# m1_18926_16202# vss nfet$197
Xnfet$214_0 m1_4620_20152# m1_4620_20152# m1_2590_19404# m1_2590_19404# m1_3454_20470#
+ vss nfet$214
Xpfet$206_1 vdd m1_n4485_21904# vdd m1_9624_19404# pfet$206
Xnfet$221_1 m1_n8625_26174# vss m1_n7082_23622# vss nfet$221
Xnfet$193_27 m1_12875_24346# m1_12875_24346# vss vss m1_12357_24542# vss nfet$193
Xnfet$193_16 m1_24808_24224# m1_24808_24224# m1_24452_24542# m1_24452_24542# m1_24906_24542#
+ vss nfet$193
Xpfet$181_99 vdd vdd m1_26705_24542# m1_24309_25858# pfet$181
Xnfet$202_12 m1_32675_25947# vss m1_28624_21786# vss nfet$202
Xpfet$181_88 vdd vdd m1_28634_25662# m1_28492_25858# pfet$181
Xpfet$181_77 vdd vdd m1_20269_24542# m1_20625_24224# pfet$181
Xpfet$181_66 vdd vdd m1_15461_25858# m1_11039_21786# pfet$181
Xpfet$181_55 vdd m1_24451_25662# m1_24188_23922# m1_23964_25662# pfet$181
Xpfet$181_44 vdd m1_15943_25858# vdd m1_17546_25658# pfet$181
Xpfet$181_33 vdd vdd m1_7522_21786# m1_7577_25858# pfet$181
Xpfet$181_22 vdd vdd m1_3537_24542# m1_3893_24224# pfet$181
Xpfet$181_11 vdd vdd m1_7719_25662# m1_7577_25858# pfet$181
Xnfet$194_81 m1_n7513_20152# vss m1_25424_24346# vss nfet$194
Xnfet$194_70 m1_21590_21786# vss m1_28010_25858# vss nfet$194
Xnfet$213_22 m1_15564_15778# m1_15564_15778# m1_15454_18030# m1_15454_18030# m1_15690_17358#
+ vss nfet$213
Xnfet$213_11 m1_6377_16202# m1_6377_16202# vss vss m1_5859_16398# vss nfet$213
Xnfet$199_15 m1_17697_15478# vss m1_22205_20152# vss nfet$199
Xnfet$198_6 m1_5771_21786# vss m1_5901_21590# vss nfet$198
Xpfet$187_10 vdd vdd m1_29239_20152# m1_26063_15478# pfet$187
Xnfet$196_3 m1_4832_17714# m1_4832_17714# vss vss m1_10488_20470# vss nfet$196
Xnfet$196_16 m1_23486_19550# m1_23486_19550# vss vss m1_23924_20470# vss nfet$196
Xnfet$216_4 m1_27031_17343# m1_27292_16202# m1_26807_17518# vss nfet$216
Xnfet$223_5 m1_n4464_25980# m1_n3541_23922# m1_n4362_24346# vss nfet$223
Xnfet$194_0 m1_3394_25858# vss m1_5790_24542# vss nfet$194
Xpfet$184_33 vdd m1_n3206_20274# m1_n3206_20274# m1_24560_19550# m1_21564_17714# m1_21564_17714#
+ pfet$184
Xpfet$184_22 vdd vdd vdd m1_14009_19550# m1_9331_15478# m1_9331_15478# pfet$184
Xpfet$184_11 vdd vdd vdd m1_10492_19550# m1_5148_15478# m1_5148_15478# pfet$184
Xpfet$186_1 vdd vdd m1_n4377_15778# m1_n7247_17714# pfet$186
Xnfet$221_11 m1_n10452_25858# vss m1_n4847_25662# vss nfet$221
Xpfet$193_2 vdd m1_n290_24224# m1_814_25658# m1_n1271_25858# pfet$193
Xnfet$197_81 m1_13198_17714# vss m1_10299_17343# vss nfet$197
Xnfet$197_70 m1_n7513_20152# vss m1_18310_16080# vss nfet$197
Xnfet$207_0 m1_21456_22513# m1_21456_22513# m1_30256_19792# m1_30256_19792# m1_30492_20470#
+ vss nfet$207
Xnfet$214_1 m1_1103_20152# m1_1103_20152# m1_n927_19404# m1_n927_19404# m1_n63_20470#
+ vss nfet$214
Xpfet$206_2 vdd m1_n5227_21418# vdd m1_2590_19404# pfet$206
Xnfet$221_2 vss vss m1_n9336_24346# vss nfet$221
Xnfet$193_17 m1_20625_24224# m1_20625_24224# m1_20269_24542# m1_20269_24542# m1_20723_24542#
+ vss nfet$193
Xnfet$202_13 m1_32675_25947# vss m1_32817_25662# vss nfet$202
Xpfet$181_89 vdd vdd m1_19839_21786# pd7 pfet$181
Xpfet$181_78 vdd m1_20269_24542# vdd m1_21241_24346# pfet$181
Xpfet$181_67 vdd m1_15822_23922# m1_16086_24542# m1_15461_25858# pfet$181
Xpfet$181_56 vdd m1_24808_24224# m1_25912_25658# m1_23827_25858# pfet$181
Xpfet$181_45 vdd vdd m1_16442_24224# m1_15822_23922# pfet$181
Xpfet$181_34 vdd m1_9180_25658# m1_9973_24542# m1_7232_25662# pfet$181
Xpfet$181_23 vdd m1_3537_24542# vdd m1_4509_24346# pfet$181
Xpfet$181_12 vdd m1_7577_25858# vdd m1_9180_25658# pfet$181
Xpfet$211_0 vdd vdd m1_n5227_20152# m1_n2543_20130# pfet$211
Xnfet$194_82 m1_11415_25662# m1_12259_24224# m1_13363_25658# vss nfet$194
Xnfet$194_71 m1_28147_25662# m1_28371_23922# m1_28635_24542# vss nfet$194
Xnfet$194_60 pd6 vss m1_16322_21786# vss nfet$194
Xnfet$213_23 m1_18926_16202# m1_18926_16202# vss vss m1_18408_16398# vss nfet$213
Xnfet$213_12 m1_n1168_15778# m1_n1168_15778# m1_n1278_18030# m1_n1278_18030# m1_n1042_17358#
+ vss nfet$213
Xnfet$199_16 m1_17381_17714# vss m1_19969_19550# vss nfet$199
Xnfet$198_7 m1_4005_21786# vss m1_4637_21786# vss nfet$198
Xpfet$187_11 vdd vdd m1_18688_20152# m1_13514_15478# pfet$187
Xnfet$196_4 m1_9418_19550# m1_9418_19550# vss vss m1_9856_20470# vss nfet$196
Xnfet$196_17 m1_12935_19550# m1_12935_19550# vss vss m1_13373_20470# vss nfet$196
Xnfet$216_5 m1_27031_17343# m1_29087_15778# m1_28470_16080# vss nfet$216
Xnfet$223_6 m1_n4464_25980# m1_n3184_24224# m1_n3651_26174# vss nfet$223
Xpfet$193_3 vdd m1_814_25658# m1_1607_24542# m1_n1134_25662# pfet$193
Xpfet$186_2 vdd vdd m1_n5351_15778# m1_n4994_16080# pfet$186
Xnfet$194_1 m1_2912_25858# m1_4997_25658# m1_5790_24542# vss nfet$194
Xpfet$184_34 vdd m1_n3206_20274# m1_n3206_20274# m1_23924_19850# m1_23486_19550# m1_23486_19550#
+ pfet$184
Xpfet$184_23 vdd vdd vdd m1_16890_19850# m1_18688_20152# m1_18688_20152# pfet$184
Xpfet$184_12 vdd m1_6107_19404# m1_6107_19404# m1_6975_19550# m1_649_17714# m1_649_17714#
+ pfet$184
Xnfet$221_12 m1_n10452_25858# vss m1_n5571_25662# vss nfet$221
Xnfet$207_1 m1_14422_22513# m1_14422_22513# m1_31535_19792# m1_31535_19792# m1_31771_20470#
+ vss nfet$207
Xnfet$214_2 m1_n3218_15478# m1_n3218_15478# m1_2590_19404# m1_2590_19404# m1_2822_20470#
+ vss nfet$214
Xnfet$221_3 fin vss m1_n10933_25858# vss nfet$221
Xnfet$197_82 m1_10299_17343# vss m1_10458_17836# vss nfet$197
Xpfet$191_0 vdd vdd vdd m1_33050_22344# m1_31535_22102# m1_31535_22102# pfet$191
Xnfet$197_71 m1_14641_17836# m1_15921_16080# m1_15454_18030# vss nfet$197
Xnfet$197_60 m1_18665_17343# vss m1_18824_17836# vss nfet$197
Xpfet$206_3 vdd vdd m1_n5227_21418# m1_6107_19404# pfet$206
Xnfet$193_18 m1_21241_24346# m1_21241_24346# vss vss m1_20723_24542# vss nfet$193
Xpfet$181_79 vdd m1_17546_25658# m1_18339_24542# m1_15598_25662# pfet$181
Xpfet$181_68 vdd vdd m1_16086_24542# m1_16442_24224# pfet$181
Xpfet$181_57 vdd vdd m1_24451_25662# m1_24309_25858# pfet$181
Xpfet$181_46 vdd m1_16442_24224# m1_17546_25658# m1_15461_25858# pfet$181
Xpfet$181_35 vdd m1_7720_24542# vdd m1_8692_24346# pfet$181
Xpfet$181_24 vdd vdd m1_5790_24542# m1_3394_25858# pfet$181
Xpfet$181_13 vdd vdd m1_12259_24224# m1_11639_23922# pfet$181
Xpfet$211_1 vdd m1_n4485_20152# vdd m1_n3206_20274# pfet$211
Xpfet$204_0 vdd vdd m1_n7320_25516# m1_n7186_25858# pfet$204
Xnfet$194_72 m1_23827_25858# m1_25912_25658# m1_26705_24542# vss nfet$194
Xnfet$194_61 m1_23964_25662# m1_24808_24224# m1_25912_25658# vss nfet$194
Xnfet$194_50 m1_n7513_20152# vss m1_21241_24346# vss nfet$194
Xnfet$213_24 m1_18310_16080# m1_18310_16080# m1_17851_17714# m1_17851_17714# m1_18408_16398#
+ vss nfet$213
Xnfet$213_13 m1_n2605_16080# m1_n2605_16080# vss vss m1_n1042_17358# vss nfet$213
Xnfet$199_17 m1_21880_15478# vss m1_25722_20152# vss nfet$199
Xnfet$198_8 m1_2254_21786# vss m1_2384_21590# vss nfet$198
Xpfet$187_12 vdd vdd m1_15171_20152# m1_9331_15478# pfet$187
Xnfet$196_5 m1_649_17714# m1_649_17714# vss vss m1_6971_20470# vss nfet$196
Xnfet$223_7 m1_n4623_25487# m1_n4362_24346# m1_n4847_25662# vss nfet$223
Xpfet$193_4 vdd m1_33174_24224# m1_34278_25658# m1_32193_25858# pfet$193
Xnfet$216_6 m1_27190_17836# m1_28113_15778# m1_27292_16202# vss nfet$216
Xnfet$194_2 m1_n7513_20152# vss m1_4509_24346# vss nfet$194
Xpfet$184_35 vdd m1_n3822_21786# m1_n3822_21786# m1_13373_19850# m1_12935_19550# m1_12935_19550#
+ pfet$184
Xpfet$184_24 vdd m1_n1927_20274# m1_n1927_20274# m1_16890_19850# m1_16452_19550# m1_16452_19550#
+ pfet$184
Xpfet$184_13 vdd m1_n927_19404# m1_n927_19404# m1_n695_19850# m1_n1133_19550# m1_n1133_19550#
+ pfet$184
Xpfet$186_3 vdd vdd m1_n6657_17518# m1_n7247_17714# pfet$186
Xnfet$221_13 fin vss m1_n4623_25487# vss nfet$221
Xnfet$207_2 m1_17939_22513# m1_17939_22513# vss vss m1_31771_20470# vss nfet$207
Xnfet$214_3 m1_8137_20152# m1_8137_20152# m1_6107_19404# m1_6107_19404# m1_6971_20470#
+ vss nfet$214
Xnfet$221_4 m1_n10572_23922# vss m1_n9952_24224# vss nfet$221
Xnfet$197_72 m1_17851_17714# vss m1_18441_17518# vss nfet$197
Xnfet$197_61 m1_20104_16080# vss m1_19747_15778# vss nfet$197
Xnfet$197_50 m1_25747_17714# vss m1_22848_17343# vss nfet$197
Xpfet$184_0 vdd m1_2590_19404# m1_2590_19404# m1_3458_19550# m1_n3534_17714# m1_n3534_17714#
+ pfet$184
Xpfet$206_4 vdd vdd m1_n4485_21904# m1_n3822_21786# pfet$206
Xnfet$193_19 m1_21729_25658# m1_21729_25658# vss vss m1_22188_25502# vss nfet$193
Xnfet$212_0 fout vss m1_35837_22102# vss nfet$212
Xpfet$181_14 vdd vdd m1_11902_25662# m1_11760_25858# pfet$181
Xpfet$211_2 vdd m1_n5227_20152# vdd m1_n1927_20274# pfet$211
Xpfet$181_69 vdd vdd m1_12875_24346# m1_n7513_20152# pfet$181
Xpfet$181_58 vdd vdd m1_23964_25662# m1_23827_25858# pfet$181
Xpfet$181_47 vdd vdd m1_15943_25858# m1_17058_24346# pfet$181
Xpfet$181_36 vdd vdd m1_8692_24346# m1_n7513_20152# pfet$181
Xpfet$181_25 vdd vdd m1_4005_21786# m1_3394_25858# pfet$181
Xpfet$204_1 vdd vdd m1_n6111_25858# m1_n6856_24542# pfet$204
Xnfet$194_73 m1_24309_25858# vss m1_21590_21786# vss nfet$194
Xnfet$194_62 m1_24188_23922# vss m1_24808_24224# vss nfet$194
Xnfet$194_51 m1_19644_25858# m1_21729_25658# m1_22522_24542# vss nfet$194
Xnfet$194_40 m1_15598_25662# m1_16442_24224# m1_17546_25658# vss nfet$194
Xnfet$213_25 m1_14743_16202# m1_14743_16202# vss vss m1_14225_16398# vss nfet$213
Xnfet$213_14 m1_n2605_16080# m1_n2605_16080# m1_n3064_17714# m1_n3064_17714# m1_n2507_16398#
+ vss nfet$213
Xnfet$198_9 m1_23356_21786# vss m1_23486_21590# vss nfet$198
Xpfet$182_90 vdd m1_19747_15778# m1_18926_16202# m1_18665_17343# pfet$182
Xpfet$187_13 vdd vdd m1_16452_19550# m1_13198_17714# pfet$187
Xnfet$196_6 m1_n1133_19550# m1_n1133_19550# vss vss m1_n695_20470# vss nfet$196
Xnfet$216_7 m1_27190_17836# m1_28470_16080# m1_28003_18030# vss nfet$216
Xnfet$194_3 m1_488_21786# vss m1_2912_25858# vss nfet$194
Xpfet$193_5 vdd m1_32817_25662# m1_32554_23922# m1_32330_25662# pfet$193
Xpfet$184_25 vdd vdd vdd m1_17526_19550# m1_13514_15478# m1_13514_15478# pfet$184
Xpfet$184_14 vdd m1_n927_19404# m1_n927_19404# m1_n59_19550# m1_n7383_17599# m1_n7383_17599#
+ pfet$184
Xpfet$186_4 vdd vdd m1_n6433_17343# m1_n3534_17714# pfet$186
Xnfet$207_3 m1_24973_22513# m1_24973_22513# vss vss m1_30492_20470# vss nfet$207
Xnfet$214_4 m1_965_15478# m1_965_15478# m1_6107_19404# m1_6107_19404# m1_6339_20470#
+ vss nfet$214
Xnfet$221_5 m1_n10933_25858# vss m1_n10796_25662# vss nfet$221
Xnfet$197_73 m1_13668_17714# vss m1_16538_15778# vss nfet$197
Xnfet$197_62 m1_18665_17343# m1_20721_15778# m1_20104_16080# vss nfet$197
Xnfet$197_51 m1_n7513_20152# vss m1_22493_16080# vss nfet$197
Xpfet$184_1 vdd vdd vdd m1_2822_19850# m1_4620_20152# m1_4620_20152# pfet$184
Xnfet$197_40 m1_n2250_17343# m1_n194_15778# m1_n811_16080# vss nfet$197
Xpfet$206_5 vdd m1_n6839_21786# vdd m1_n5764_21786# pfet$206
Xnfet$212_1 define m1_35837_22102# vss vss nfet$212
Xnfet$205_0 m1_n290_24224# m1_n290_24224# m1_n646_24542# m1_n646_24542# m1_n192_24542#
+ vss nfet$205
Xpfet$181_59 vdd vdd m1_16322_21786# pd6 pfet$181
Xpfet$181_48 vdd m1_16085_25662# m1_15822_23922# m1_15598_25662# pfet$181
Xpfet$181_37 vdd vdd m1_9973_24542# m1_7577_25858# pfet$181
Xpfet$181_26 vdd m1_4997_25658# m1_5790_24542# m1_3049_25662# pfet$181
Xpfet$181_15 vdd m1_11902_25662# m1_11639_23922# m1_11415_25662# pfet$181
Xpfet$211_3 vdd m1_n6839_20152# vdd m1_n927_19404# pfet$211
Xnfet$194_74 pd8 vss m1_23356_21786# vss nfet$194
Xnfet$194_63 m1_14556_21786# vss m1_19644_25858# vss nfet$194
Xnfet$194_52 m1_20126_25858# vss m1_22522_24542# vss nfet$194
Xnfet$194_41 pd5 vss m1_12805_21786# vss nfet$194
Xnfet$194_30 m1_n7513_20152# vss m1_17058_24346# vss nfet$194
Xnfet$213_26 m1_14127_16080# m1_14127_16080# m1_13668_17714# m1_13668_17714# m1_14225_16398#
+ vss nfet$213
Xnfet$213_15 m1_n1989_16202# m1_n1989_16202# vss vss m1_n2507_16398# vss nfet$213
Xpfet$182_91 vdd m1_24287_16080# m1_23820_18030# m1_22848_17343# pfet$182
Xpfet$182_80 vdd vdd m1_15564_15778# m1_15921_16080# pfet$182
Xpfet$187_14 vdd vdd m1_23486_19550# m1_21564_17714# pfet$187
Xnfet$196_7 m1_n7383_17599# m1_n7383_17599# vss vss m1_n63_20470# vss nfet$196
Xnfet$194_4 m1_2912_25858# vss m1_3049_25662# vss nfet$194
Xpfet$193_6 vdd m1_34278_25658# m1_35071_24542# m1_32330_25662# pfet$193
Xpfet$184_26 vdd m1_n1927_20274# m1_n1927_20274# m1_17526_19550# m1_13198_17714# m1_13198_17714#
+ pfet$184
Xpfet$184_15 vdd vdd vdd m1_n59_19550# m1_n7401_15478# m1_n7401_15478# pfet$184
Xpfet$186_5 vdd vdd m1_n6788_16080# m1_n7513_20152# pfet$186
Xnfet$221_6 m1_n10452_25858# vss m1_n10309_25662# vss nfet$221
Xnfet$197_74 m1_14482_17343# vss m1_14641_17836# vss nfet$197
Xnfet$197_63 m1_13668_17714# vss m1_14258_17518# vss nfet$197
Xnfet$197_52 m1_23007_17836# m1_24287_16080# m1_23820_18030# vss nfet$197
Xnfet$207_4 m1_32818_20470# m1_32818_20470# vss vss m1_34329_20470# vss nfet$207
Xnfet$214_5 m1_5148_15478# m1_5148_15478# m1_9624_19404# m1_9624_19404# m1_9856_20470#
+ vss nfet$214
Xnfet$197_30 sd6 vss m1_5148_15478# vss nfet$197
Xnfet$197_41 m1_n2091_17836# m1_n1168_15778# m1_n1989_16202# vss nfet$197
Xpfet$206_6 vdd vdd m1_n6973_21481# m1_n6839_21786# pfet$206
Xpfet$184_2 vdd m1_2590_19404# m1_2590_19404# m1_2822_19850# m1_2384_19550# m1_2384_19550#
+ pfet$184
Xnfet$205_1 m1_814_25658# m1_814_25658# vss vss m1_1273_25502# vss nfet$205
Xpfet$181_49 vdd m1_20126_25858# vdd m1_21729_25658# pfet$181
Xpfet$181_38 vdd vdd m1_16085_25662# m1_15943_25858# pfet$181
Xpfet$181_27 vdd vdd m1_11278_25858# m1_7522_21786# pfet$181
Xpfet$181_16 vdd vdd m1_5771_21786# pd3 pfet$181
Xpfet$211_4 vdd vdd m1_n6839_20152# m1_n6973_21481# pfet$211
Xnfet$194_75 m1_28371_23922# vss m1_28991_24224# vss nfet$194
Xnfet$194_64 m1_19644_25858# vss m1_19781_25662# vss nfet$194
Xnfet$194_53 m1_23827_25858# m1_24451_25662# m1_24188_23922# vss nfet$194
Xnfet$194_42 m1_15943_25858# vss m1_16085_25662# vss nfet$194
Xnfet$194_31 m1_15943_25858# vss m1_18339_24542# vss nfet$194
Xnfet$213_27 m1_18310_16080# m1_18310_16080# vss vss m1_19873_17358# vss nfet$213
Xnfet$213_16 m1_19747_15778# m1_19747_15778# m1_19637_18030# m1_19637_18030# m1_19873_17358#
+ vss nfet$213
Xnfet$194_20 pd3 vss m1_5771_21786# vss nfet$194
Xpfet$182_81 vdd vdd m1_13668_17714# m1_14127_16080# pfet$182
Xpfet$182_70 vdd vdd m1_18824_17836# m1_18665_17343# pfet$182
Xpfet$202_0 vdd vdd vdd m1_n6624_23622# m1_n7082_23622# m1_n7082_23622# pfet$202
Xpfet$182_92 vdd m1_15454_18030# vdd m1_14127_16080# pfet$182
Xpfet$187_15 vdd vdd m1_22205_20152# m1_17697_15478# pfet$187
Xnfet$196_8 m1_27003_19550# m1_27003_19550# vss vss m1_27441_20470# vss nfet$196
Xnfet$194_5 m1_2912_25858# m1_3536_25662# m1_3273_23922# vss nfet$194
Xpfet$193_7 vdd m1_32554_23922# m1_32818_24542# m1_32193_25858# pfet$193
Xpfet$184_27 vdd vdd vdd m1_20407_19850# m1_22205_20152# m1_22205_20152# pfet$184
Xpfet$184_16 vdd vdd vdd m1_28077_19550# m1_26063_15478# m1_26063_15478# pfet$184
Xnfet$228_0 m1_n4485_20152# m1_n6380_21786# vss vss nfet$228
Xpfet$186_6 vdd vdd m1_n7383_17599# m1_n7247_17714# pfet$186
Xpfet$207_10 vdd vdd m1_n10933_25858# fin pfet$207
Xnfet$197_75 sd3 vss m1_17697_15478# vss nfet$197
Xnfet$197_64 m1_13668_17714# vss m1_13198_17714# vss nfet$197
Xnfet$197_53 m1_22848_17343# vss m1_23007_17836# vss nfet$197
Xnfet$207_5 m1_32818_21586# m1_32818_21586# m1_34093_19792# m1_34093_19792# m1_34329_20470#
+ vss nfet$207
Xnfet$197_31 m1_1933_17343# m1_3989_15778# m1_3372_16080# vss nfet$197
Xnfet$197_20 m1_1119_17714# vss m1_1709_17518# vss nfet$197
Xnfet$214_6 m1_11654_20152# m1_11654_20152# m1_9624_19404# m1_9624_19404# m1_10488_20470#
+ vss nfet$214
Xnfet$197_42 m1_n811_16080# vss m1_n1168_15778# vss nfet$197
Xnfet$221_7 m1_n7320_25516# vss m1_n2567_23922# vss nfet$221
Xpfet$206_7 vdd vdd m1_n6839_21786# m1_n6380_21786# pfet$206
Xpfet$184_3 vdd vdd vdd m1_3458_19550# m1_n3218_15478# m1_n3218_15478# pfet$184
Xnfet$205_2 m1_326_24346# m1_326_24346# m1_n789_25858# m1_n789_25858# m1_1273_25502#
+ vss nfet$205
Xpfet$181_39 vdd vdd m1_15598_25662# m1_15461_25858# pfet$181
Xpfet$181_28 vdd m1_11639_23922# m1_11903_24542# m1_11278_25858# pfet$181
Xpfet$181_17 vdd vdd m1_7577_25858# m1_8692_24346# pfet$181
Xpfet$182_0 vdd vdd m1_12355_15778# m1_9485_17714# pfet$182
Xnfet$194_76 m1_28492_25858# vss m1_28634_25662# vss nfet$194
Xnfet$194_65 m1_28492_25858# vss m1_25107_21786# vss nfet$194
Xnfet$194_54 m1_24309_25858# vss m1_24451_25662# vss nfet$194
Xnfet$194_43 m1_15461_25858# vss m1_15598_25662# vss nfet$194
Xnfet$194_32 m1_15461_25858# m1_17546_25658# m1_18339_24542# vss nfet$194
Xnfet$213_17 m1_22493_16080# m1_22493_16080# vss vss m1_24056_17358# vss nfet$213
Xnfet$210_0 m1_34093_19792# vss m1_34843_21786# vss nfet$210
Xnfet$194_21 m1_11278_25858# m1_11902_25662# m1_11639_23922# vss nfet$194
Xnfet$194_10 m1_7577_25858# vss m1_9973_24542# vss nfet$194
Xpfet$202_1 vdd m1_n6856_24542# m1_n6856_24542# m1_n6624_23622# m1_n8283_19850# m1_n8283_19850#
+ pfet$202
Xpfet$182_93 vdd m1_23820_18030# vdd m1_22493_16080# pfet$182
Xpfet$182_82 vdd m1_13668_17714# vdd m1_14743_16202# pfet$182
Xpfet$182_71 vdd vdd m1_19747_15778# m1_20104_16080# pfet$182
Xpfet$182_60 vdd vdd m1_n194_15778# m1_n3064_17714# pfet$182
Xpfet$187_16 vdd vdd m1_19969_19550# m1_17381_17714# pfet$187
Xnfet$196_9 m1_25747_17714# m1_25747_17714# vss vss m1_28073_20470# vss nfet$196
Xpfet$186_7 vdd vdd m1_27190_17836# m1_27031_17343# pfet$186
Xnfet$194_6 m1_3049_25662# m1_3893_24224# m1_4997_25658# vss nfet$194
Xnfet$228_1 m1_n5227_20152# vss m1_n6380_21786# vss nfet$228
Xpfet$207_11 vdd vdd m1_n9336_24346# vss pfet$207
Xpfet$184_28 vdd vdd vdd m1_21043_19550# m1_17697_15478# m1_17697_15478# pfet$184
Xpfet$184_17 vdd m1_n3822_20130# m1_n3822_20130# m1_28077_19550# m1_25747_17714# m1_25747_17714#
+ pfet$184
Xnfet$207_6 m1_354_22513# m1_354_22513# m1_31535_22102# m1_31535_22102# m1_31771_21430#
+ vss nfet$207
Xnfet$214_7 m1_n7401_15478# m1_n7401_15478# m1_n927_19404# m1_n927_19404# m1_n695_20470#
+ vss nfet$214
Xnfet$197_10 m1_11738_16080# vss m1_11381_15778# vss nfet$197
Xnfet$221_8 m1_n4623_25487# vss m1_n4464_25980# vss nfet$221
Xnfet$197_76 m1_14482_17343# m1_16538_15778# m1_15921_16080# vss nfet$197
Xnfet$197_65 m1_14482_17343# m1_14743_16202# m1_14258_17518# vss nfet$197
Xnfet$197_54 m1_22848_17343# m1_23109_16202# m1_22624_17518# vss nfet$197
Xpfet$184_4 vdd m1_6107_19404# m1_6107_19404# m1_6339_19850# m1_5901_19550# m1_5901_19550#
+ pfet$184
Xnfet$197_32 m1_2092_17836# m1_3015_15778# m1_2194_16202# vss nfet$197
Xnfet$197_21 m1_1933_17343# m1_2194_16202# m1_1709_17518# vss nfet$197
Xnfet$197_43 sd8 vss m1_n3218_15478# vss nfet$197
Xnfet$205_3 m1_326_24346# m1_326_24346# vss vss m1_n192_24542# vss nfet$205
Xpfet$181_29 vdd vdd m1_11903_24542# m1_12259_24224# pfet$181
Xpfet$181_18 vdd vdd m1_11415_25662# m1_11278_25858# pfet$181
Xpfet$182_1 vdd vdd m1_11381_15778# m1_11738_16080# pfet$182
Xnfet$194_77 m1_28010_25858# vss m1_28147_25662# vss nfet$194
Xnfet$194_66 m1_28010_25858# m1_30095_25658# m1_30888_24542# vss nfet$194
Xnfet$194_55 m1_23827_25858# vss m1_23964_25662# vss nfet$194
Xnfet$194_44 m1_15822_23922# vss m1_16442_24224# vss nfet$194
Xnfet$194_33 m1_11760_25858# vss m1_14156_24542# vss nfet$194
Xnfet$210_1 m1_30256_19792# vss m1_32818_20470# vss nfet$210
Xnfet$194_22 m1_11760_25858# vss m1_11902_25662# vss nfet$194
Xnfet$194_11 m1_7522_21786# vss m1_11278_25858# vss nfet$194
Xnfet$203_0 m1_n1134_25662# m1_n910_23922# m1_n646_24542# vss nfet$203
Xnfet$213_18 m1_23930_15778# m1_23930_15778# m1_23820_18030# m1_23820_18030# m1_24056_17358#
+ vss nfet$213
Xpfet$182_94 vdd vdd m1_22624_17518# m1_22034_17714# pfet$182
Xpfet$182_83 vdd m1_16538_15778# m1_15921_16080# m1_14641_17836# pfet$182
Xpfet$182_72 vdd m1_20721_15778# m1_20104_16080# m1_18824_17836# pfet$182
Xpfet$182_61 vdd m1_n811_16080# m1_n1278_18030# m1_n2250_17343# pfet$182
Xpfet$182_50 vdd m1_n1168_15778# m1_n1989_16202# m1_n2250_17343# pfet$182
Xpfet$187_17 vdd vdd m1_25722_20152# m1_21880_15478# pfet$187
Xnfet$194_7 m1_3049_25662# m1_3273_23922# m1_3537_24542# vss nfet$194
Xpfet$207_12 vdd vdd m1_n7082_23622# m1_n8625_26174# pfet$207
Xpfet$184_29 vdd vdd vdd m1_23924_19850# m1_25722_20152# m1_25722_20152# pfet$184
Xpfet$184_18 vdd vdd vdd m1_27441_19850# m1_29239_20152# m1_29239_20152# pfet$184
Xpfet$186_8 vdd vdd m1_28113_15778# m1_28470_16080# pfet$186
Xnfet$207_7 m1_3871_22513# m1_3871_22513# vss vss m1_31771_21430# vss nfet$207
Xnfet$214_8 m1_26063_15478# m1_26063_15478# m1_n3822_20130# m1_n3822_20130# m1_27441_20470#
+ vss nfet$214
Xnfet$221_9 m1_n3184_24224# vss m1_n3541_23922# vss nfet$221
Xnfet$197_77 sd4 vss m1_13514_15478# vss nfet$197
Xnfet$197_66 m1_n7513_20152# vss m1_14127_16080# vss nfet$197
Xnfet$197_55 m1_22034_17714# vss m1_24904_15778# vss nfet$197
Xnfet$197_44 m1_n2091_17836# m1_n811_16080# m1_n1278_18030# vss nfet$197
Xpfet$184_5 vdd vdd vdd m1_n695_19850# m1_1103_20152# m1_1103_20152# pfet$184
Xnfet$197_33 sd7 vss m1_965_15478# vss nfet$197
Xnfet$197_22 m1_6116_17343# m1_6377_16202# m1_5892_17518# vss nfet$197
Xnfet$197_11 m1_10299_17343# m1_12355_15778# m1_11738_16080# vss nfet$197
Xnfet$205_4 m1_33174_24224# m1_33174_24224# m1_32818_24542# m1_32818_24542# m1_33272_24542#
+ vss nfet$205
Xpfet$181_19 vdd vdd m1_7095_25858# m1_4005_21786# pfet$181
Xpfet$182_2 vdd m1_12355_15778# m1_11738_16080# m1_10458_17836# pfet$182
Xnfet$194_78 m1_28010_25858# m1_28634_25662# m1_28371_23922# vss nfet$194
Xnfet$194_67 m1_28492_25858# vss m1_30888_24542# vss nfet$194
Xnfet$194_56 m1_19781_25662# m1_20625_24224# m1_21729_25658# vss nfet$194
Xnfet$194_45 m1_15461_25858# m1_16085_25662# m1_15822_23922# vss nfet$194
Xnfet$194_34 m1_11278_25858# m1_13363_25658# m1_14156_24542# vss nfet$194
Xnfet$210_2 m1_31535_19792# m1_32818_20470# vss vss nfet$210
Xnfet$194_23 m1_11278_25858# vss m1_11415_25662# vss nfet$194
Xnfet$194_12 m1_7577_25858# vss m1_7522_21786# vss nfet$194
Xnfet$213_19 m1_23109_16202# m1_23109_16202# vss vss m1_22591_16398# vss nfet$213
Xnfet$203_1 m1_n1271_25858# m1_n647_25662# m1_n910_23922# vss nfet$203
Xpfet$182_95 vdd vdd m1_21564_17714# m1_22034_17714# pfet$182
Xpfet$182_84 vdd vdd m1_17381_17714# m1_17851_17714# pfet$182
Xpfet$182_73 vdd vdd m1_16538_15778# m1_13668_17714# pfet$182
Xpfet$182_62 vdd vdd m1_23007_17836# m1_22848_17343# pfet$182
Xpfet$182_40 vdd m1_10560_16202# m1_10075_17518# m1_10458_17836# pfet$182
Xpfet$182_51 vdd vdd m1_n1168_15778# m1_n811_16080# pfet$182
Xpfet$200_0 vdd m1_n4377_15778# m1_n4994_16080# m1_n6274_17836# pfet$200
Xnfet$194_8 m1_3394_25858# vss m1_3536_25662# vss nfet$194
Xpfet$207_13 vdd vdd m1_n8055_24542# m1_n8625_26174# pfet$207
Xpfet$184_19 vdd m1_n3822_20130# m1_n3822_20130# m1_27441_19850# m1_27003_19550# m1_27003_19550#
+ pfet$184
Xpfet$186_9 vdd vdd m1_29087_15778# m1_26217_17714# pfet$186
Xpfet$198_0 vdd m1_32818_20470# m1_32818_20470# m1_33050_19550# m1_30256_19792# m1_30256_19792#
+ pfet$198
Xnfet$214_9 m1_29239_20152# m1_29239_20152# m1_n3822_20130# m1_n3822_20130# m1_28073_20470#
+ vss nfet$214
Xnfet$197_78 m1_14641_17836# m1_15564_15778# m1_14743_16202# vss nfet$197
Xnfet$197_67 m1_17381_17714# vss m1_14482_17343# vss nfet$197
Xnfet$197_56 m1_24287_16080# vss m1_23930_15778# vss nfet$197
Xnfet$197_45 m1_n3064_17714# vss m1_n194_15778# vss nfet$197
Xnfet$197_34 m1_n2250_17343# vss m1_n2091_17836# vss nfet$197
Xnfet$197_23 m1_5302_17714# vss m1_4832_17714# vss nfet$197
Xnfet$197_12 m1_9485_17714# vss m1_12355_15778# vss nfet$197
Xpfet$184_6 vdd vdd vdd m1_6339_19850# m1_8137_20152# m1_8137_20152# pfet$184
Xnfet$226_0 m1_n4485_21904# m1_n5764_21786# vss vss nfet$226
Xnfet$205_5 m1_33790_24346# m1_33790_24346# vss vss m1_33272_24542# vss nfet$205
Xpfet$182_3 vdd m1_11381_15778# m1_10560_16202# m1_10299_17343# pfet$182
Xnfet$194_79 pd7 vss m1_19839_21786# vss nfet$194
Xnfet$194_68 m1_n7513_20152# vss m1_29607_24346# vss nfet$194
Xnfet$210_3 m1_30256_22102# vss m1_32818_21586# vss nfet$210
Xnfet$194_57 m1_20126_25858# vss m1_20268_25662# vss nfet$194
Xnfet$194_46 m1_20126_25858# vss m1_18073_21786# vss nfet$194
Xnfet$194_35 m1_15598_25662# m1_15822_23922# m1_16086_24542# vss nfet$194
Xnfet$194_24 m1_7095_25858# m1_7719_25662# m1_7456_23922# vss nfet$194
Xnfet$194_13 m1_11415_25662# m1_11639_23922# m1_11903_24542# vss nfet$194
Xnfet$203_2 m1_n1271_25858# m1_814_25658# m1_1607_24542# vss nfet$203
Xpfet$182_96 vdd vdd m1_18665_17343# m1_21564_17714# pfet$182
Xpfet$182_85 vdd m1_18926_16202# m1_18441_17518# m1_18824_17836# pfet$182
Xpfet$182_74 vdd vdd m1_14641_17836# m1_14482_17343# pfet$182
Xpfet$182_63 vdd m1_23930_15778# m1_23109_16202# m1_22848_17343# pfet$182
Xpfet$182_30 vdd vdd m1_1933_17343# m1_4832_17714# pfet$182
Xpfet$182_41 vdd vdd m1_10075_17518# m1_9485_17714# pfet$182
Xpfet$182_52 vdd m1_n3064_17714# vdd m1_n1989_16202# pfet$182
Xpfet$200_1 vdd m1_n5351_15778# m1_n6172_16202# m1_n6433_17343# pfet$200
Xnfet$194_9 m1_3273_23922# vss m1_3893_24224# vss nfet$194
Xpfet$198_1 vdd vdd vdd m1_33050_19550# m1_31535_19792# m1_31535_19792# pfet$198
Xnfet$197_79 m1_15921_16080# vss m1_15564_15778# vss nfet$197
Xnfet$197_68 m1_18665_17343# m1_18926_16202# m1_18441_17518# vss nfet$197
Xnfet$197_57 m1_22848_17343# m1_24904_15778# m1_24287_16080# vss nfet$197
Xnfet$197_46 m1_22034_17714# vss m1_21564_17714# vss nfet$197
Xnfet$197_24 m1_4832_17714# vss m1_1933_17343# vss nfet$197
Xnfet$197_13 m1_10458_17836# m1_11381_15778# m1_10560_16202# vss nfet$197
Xnfet$197_35 m1_n7513_20152# vss m1_5761_16080# vss nfet$197
Xnfet$226_1 m1_n5227_21418# vss m1_n5764_21786# vss nfet$226
Xnfet$219_0 m1_n7082_23622# m1_n6856_24542# vss vss nfet$219
Xpfet$182_110 vdd vdd m1_10458_17836# m1_10299_17343# pfet$182
Xpfet$184_7 vdd vdd vdd m1_6975_19550# m1_965_15478# m1_965_15478# pfet$184
Xnfet$205_6 m1_33790_24346# m1_33790_24346# m1_32675_25947# m1_32675_25947# m1_34737_25502#
+ vss nfet$205
Xpfet$182_4 vdd m1_9485_17714# vdd m1_10560_16202# pfet$182
Xnfet$194_69 m1_24309_25858# vss m1_26705_24542# vss nfet$194
Xnfet$194_58 m1_20005_23922# vss m1_20625_24224# vss nfet$194
Xnfet$194_47 m1_23964_25662# m1_24188_23922# m1_24452_24542# vss nfet$194
Xnfet$194_36 m1_11760_25858# vss m1_11039_21786# vss nfet$194
Xnfet$194_25 m1_7232_25662# m1_8076_24224# m1_9180_25658# vss nfet$194
Xnfet$194_14 m1_n7513_20152# vss m1_8692_24346# vss nfet$194
Xnfet$203_3 m1_n1134_25662# m1_n290_24224# m1_814_25658# vss nfet$203
Xpfet$182_97 vdd vdd m1_22493_16080# m1_n7513_20152# pfet$182
Xpfet$182_86 vdd m1_19637_18030# vdd m1_18310_16080# pfet$182
Xpfet$182_75 vdd vdd m1_17697_15478# sd3 pfet$182
Xpfet$182_64 vdd vdd m1_23930_15778# m1_24287_16080# pfet$182
Xpfet$182_20 vdd vdd m1_1119_17714# m1_1578_16080# pfet$182
Xpfet$182_31 vdd m1_3372_16080# m1_2905_18030# m1_1933_17343# pfet$182
Xpfet$182_42 vdd m1_11271_18030# vdd m1_9944_16080# pfet$182
Xpfet$182_53 vdd vdd m1_n3218_15478# sd8 pfet$182
Xnfet$201_0 m1_n3534_17714# vss m1_n6433_17343# vss nfet$201
Xpfet$200_2 vdd m1_n4994_16080# m1_n5461_18030# m1_n6433_17343# pfet$200
Xnfet$199_0 m1_n3534_17714# vss m1_2384_19550# vss nfet$199
Xpfet$198_2 vdd m1_32818_21586# m1_32818_21586# m1_33050_22344# m1_30256_22102# m1_30256_22102#
+ pfet$198
Xnfet$197_69 m1_17851_17714# vss m1_17381_17714# vss nfet$197
Xnfet$197_58 m1_23007_17836# m1_23930_15778# m1_23109_16202# vss nfet$197
Xnfet$197_47 m1_22034_17714# vss m1_22624_17518# vss nfet$197
Xnfet$197_25 m1_2092_17836# m1_3372_16080# m1_2905_18030# vss nfet$197
Xnfet$197_14 m1_6116_17343# m1_8172_15778# m1_7555_16080# vss nfet$197
Xnfet$197_36 m1_n3064_17714# vss m1_n2474_17518# vss nfet$197
Xpfet$184_8 vdd m1_9624_19404# m1_9624_19404# m1_10492_19550# m1_4832_17714# m1_4832_17714#
+ pfet$184
Xnfet$226_2 m1_n6839_21786# vss m1_n6973_21481# vss nfet$226
Xnfet$219_1 m1_n8283_19850# vss m1_n6856_24542# vss nfet$219
Xnfet$205_7 m1_34278_25658# m1_34278_25658# vss vss m1_34737_25502# vss nfet$205
Xnfet$206_10 m1_21590_21786# m1_21590_21786# vss vss m1_20428_21586# vss nfet$206
Xpfet$182_100 vdd vdd m1_23820_18030# m1_23930_15778# pfet$182
Xpfet$182_5 vdd m1_7198_15778# m1_6377_16202# m1_6116_17343# pfet$182
Xnfet$203_4 m1_32193_25858# m1_34278_25658# m1_35071_24542# vss nfet$203
Xnfet$194_59 m1_19644_25858# m1_20268_25662# m1_20005_23922# vss nfet$194
Xnfet$194_48 m1_18073_21786# vss m1_23827_25858# vss nfet$194
Xnfet$194_37 m1_11039_21786# vss m1_15461_25858# vss nfet$194
Xnfet$194_26 m1_7095_25858# m1_9180_25658# m1_9973_24542# vss nfet$194
Xnfet$194_15 m1_7232_25662# m1_7456_23922# m1_7720_24542# vss nfet$194
Xpfet$182_98 vdd m1_20104_16080# m1_19637_18030# m1_18665_17343# pfet$182
Xpfet$182_87 vdd vdd m1_18310_16080# m1_n7513_20152# pfet$182
Xpfet$182_76 vdd m1_17851_17714# vdd m1_18926_16202# pfet$182
Xpfet$182_65 vdd m1_24904_15778# m1_24287_16080# m1_23007_17836# pfet$182
Xpfet$182_21 vdd vdd m1_965_15478# sd7 pfet$182
Xpfet$182_10 vdd m1_8172_15778# m1_7555_16080# m1_6275_17836# pfet$182
Xpfet$182_32 vdd vdd m1_2905_18030# m1_3015_15778# pfet$182
Xpfet$182_43 vdd vdd m1_11271_18030# m1_11381_15778# pfet$182
Xpfet$182_54 vdd vdd m1_n1278_18030# m1_n1168_15778# pfet$182
Xnfet$201_1 m1_n7513_20152# vss m1_n6788_16080# vss nfet$201
Xpfet$200_3 vdd m1_n6172_16202# m1_n6657_17518# m1_n6274_17836# pfet$200
Xnfet$214_10 m1_9331_15478# m1_9331_15478# m1_n3822_21786# m1_n3822_21786# m1_13373_20470#
+ vss nfet$214
Xnfet$199_1 m1_n3218_15478# vss m1_4620_20152# vss nfet$199
Xnfet$197_15 m1_5302_17714# vss m1_8172_15778# vss nfet$197
Xnfet$197_59 m1_17851_17714# vss m1_20721_15778# vss nfet$197
Xnfet$197_48 m1_18824_17836# m1_20104_16080# m1_19637_18030# vss nfet$197
Xnfet$197_26 m1_5302_17714# vss m1_5892_17518# vss nfet$197
Xpfet$184_9 vdd m1_9624_19404# m1_9624_19404# m1_9856_19850# m1_9418_19550# m1_9418_19550#
+ pfet$184
Xnfet$197_37 m1_n7513_20152# vss m1_n2605_16080# vss nfet$197
Xpfet$196_0 vdd vdd vdd m1_36073_22344# define define pfet$196
Xpfet$185_10 vdd vdd m1_23486_21590# m1_23356_21786# pfet$185
Xnfet$206_11 m1_22222_21786# m1_22222_21786# vss vss m1_21060_21586# vss nfet$206
Xpfet$182_101 vdd vdd m1_19637_18030# m1_19747_15778# pfet$182
Xnfet$224_0 m1_n7186_25858# vss m1_n7320_25516# vss nfet$224
Xpfet$182_6 vdd vdd m1_7198_15778# m1_7555_16080# pfet$182
Xpfet$209_0 vdd vdd vdd m1_n8047_19550# m1_n7513_20152# m1_n7513_20152# pfet$209
Xnfet$203_5 m1_32330_25662# m1_33174_24224# m1_34278_25658# vss nfet$203
Xnfet$194_49 m1_19781_25662# m1_20005_23922# m1_20269_24542# vss nfet$194
Xnfet$194_38 m1_n7513_20152# vss m1_12875_24346# vss nfet$194
Xnfet$194_27 m1_7577_25858# vss m1_7719_25662# vss nfet$194
Xnfet$194_16 m1_4005_21786# vss m1_7095_25858# vss nfet$194
Xpfet$182_99 vdd m1_23109_16202# m1_22624_17518# m1_23007_17836# pfet$182
Xpfet$182_88 vdd vdd m1_18441_17518# m1_17851_17714# pfet$182
Xpfet$182_77 vdd vdd m1_17851_17714# m1_18310_16080# pfet$182
Xpfet$182_66 vdd vdd m1_24904_15778# m1_22034_17714# pfet$182
Xpfet$182_22 vdd vdd m1_3015_15778# m1_3372_16080# pfet$182
Xpfet$182_11 vdd vdd m1_9485_17714# m1_9944_16080# pfet$182
Xpfet$182_33 vdd vdd m1_5892_17518# m1_5302_17714# pfet$182
Xpfet$182_44 vdd vdd m1_649_17714# m1_1119_17714# pfet$182
Xpfet$182_55 vdd vdd m1_n2474_17518# m1_n3064_17714# pfet$182
Xnfet$201_2 m1_n4994_16080# vss m1_n5351_15778# vss nfet$201
Xnfet$214_11 m1_15171_20152# m1_15171_20152# m1_n3822_21786# m1_n3822_21786# m1_14005_20470#
+ vss nfet$214
Xpfet$200_4 vdd m1_28113_15778# m1_27292_16202# m1_27031_17343# pfet$200
Xnfet$199_2 m1_n7401_15478# vss m1_1103_20152# vss nfet$199
Xnfet$197_49 m1_21564_17714# vss m1_18665_17343# vss nfet$197
Xnfet$197_27 m1_1119_17714# vss m1_3989_15778# vss nfet$197
Xnfet$197_16 m1_6275_17836# m1_7198_15778# m1_6377_16202# vss nfet$197
Xnfet$197_38 m1_n2250_17343# m1_n1989_16202# m1_n2474_17518# vss nfet$197
Xpfet$196_1 vdd m1_35837_22102# m1_35837_22102# m1_36073_22344# fout fout pfet$196
Xpfet$185_11 vdd vdd m1_18705_21786# m1_18073_21786# pfet$185
Xnfet$206_12 m1_18073_21786# m1_18073_21786# vss vss m1_16911_21586# vss nfet$206
Xpfet$182_102 vdd vdd m1_13198_17714# m1_13668_17714# pfet$182
Xpfet$189_0 vdd vdd m1_n647_25662# m1_n789_25858# pfet$189
Xpfet$182_7 vdd vdd m1_6275_17836# m1_6116_17343# pfet$182
Xnfet$217_0 m1_n5351_15778# m1_n5351_15778# m1_n5461_18030# m1_n5461_18030# m1_n5225_17358#
+ vss nfet$217
Xpfet$209_1 vdd m1_n8283_19850# m1_n8283_19850# m1_n8047_19550# m1_n8283_20611# m1_n8283_20611#
+ pfet$209
Xnfet$224_1 m1_n6856_24542# vss m1_n6111_25858# vss nfet$224
Xnfet$194_39 pd4 vss m1_9288_21786# vss nfet$194
Xnfet$194_28 m1_3394_25858# vss m1_4005_21786# vss nfet$194
Xnfet$194_17 m1_11639_23922# vss m1_12259_24224# vss nfet$194
Xnfet$203_6 m1_32193_25858# m1_32817_25662# m1_32554_23922# vss nfet$203
Xpfet$182_89 vdd vdd m1_22848_17343# m1_25747_17714# pfet$182
Xpfet$182_78 vdd vdd m1_13514_15478# sd4 pfet$182
Xpfet$182_67 vdd m1_22034_17714# vdd m1_23109_16202# pfet$182
Xpfet$182_12 vdd m1_3989_15778# m1_3372_16080# m1_2092_17836# pfet$182
Xpfet$182_23 vdd m1_5302_17714# vdd m1_6377_16202# pfet$182
Xpfet$182_34 vdd vdd m1_5761_16080# m1_n7513_20152# pfet$182
Xpfet$182_45 vdd vdd m1_9944_16080# m1_n7513_20152# pfet$182
Xpfet$182_56 vdd m1_n1278_18030# vdd m1_n2605_16080# pfet$182
Xnfet$201_3 m1_n6433_17343# vss m1_n6274_17836# vss nfet$201
Xnfet$214_12 m1_18688_20152# m1_18688_20152# m1_n1927_20274# m1_n1927_20274# m1_17522_20470#
+ vss nfet$214
Xpfet$200_5 vdd m1_29087_15778# m1_28470_16080# m1_27190_17836# pfet$200
Xnfet$199_3 m1_649_17714# vss m1_5901_19550# vss nfet$199
Xnfet$197_28 m1_1933_17343# vss m1_2092_17836# vss nfet$197
Xnfet$197_17 m1_649_17714# vss m1_n2250_17343# vss nfet$197
Xnfet$197_39 m1_n3064_17714# vss m1_n3534_17714# vss nfet$197
Xpfet$185_12 vdd vdd m1_16452_21590# m1_16322_21786# pfet$185
Xnfet$206_13 m1_18705_21786# m1_18705_21786# vss vss m1_17543_21586# vss nfet$206
Xpfet$182_103 vdd m1_14743_16202# m1_14258_17518# m1_14641_17836# pfet$182
Xnfet$197_0 m1_9485_17714# vss m1_9015_17714# vss nfet$197
Xpfet$189_1 vdd vdd m1_n1134_25662# m1_n1271_25858# pfet$189
Xpfet$182_8 vdd vdd m1_9331_15478# sd5 pfet$182
Xnfet$217_1 m1_n6788_16080# m1_n6788_16080# vss vss m1_n5225_17358# vss nfet$217
Xpfet$209_2 vdd m1_n8283_20611# m1_n8283_20611# m1_n8047_22344# m1_n8145_21908# m1_n8145_21908#
+ pfet$209
Xnfet$203_7 m1_32330_25662# m1_32554_23922# m1_32818_24542# vss nfet$203
Xnfet$194_29 m1_15943_25858# vss m1_14556_21786# vss nfet$194
Xnfet$194_18 m1_7095_25858# vss m1_7232_25662# vss nfet$194
Xpfet$182_79 vdd m1_15564_15778# m1_14743_16202# m1_14482_17343# pfet$182
Xpfet$182_68 vdd vdd m1_22034_17714# m1_22493_16080# pfet$182
Xpfet$182_13 vdd vdd m1_5148_15478# sd6 pfet$182
Xpfet$182_24 vdd m1_6377_16202# m1_5892_17518# m1_6275_17836# pfet$182
Xpfet$182_35 vdd vdd m1_9015_17714# m1_9485_17714# pfet$182
Xpfet$182_46 vdd vdd m1_n2250_17343# m1_649_17714# pfet$182
Xpfet$182_57 vdd m1_n1989_16202# m1_n2474_17518# m1_n2091_17836# pfet$182
Xnfet$201_4 m1_n7247_17714# vss m1_n4377_15778# vss nfet$201
Xnfet$214_13 m1_13514_15478# m1_13514_15478# m1_n1927_20274# m1_n1927_20274# m1_16890_20470#
+ vss nfet$214
Xpfet$200_6 vdd m1_28470_16080# m1_28003_18030# m1_27031_17343# pfet$200
Xnfet$199_4 m1_4832_17714# vss m1_9418_19550# vss nfet$199
Xnfet$197_29 m1_3372_16080# vss m1_3015_15778# vss nfet$197
Xnfet$197_18 m1_1119_17714# vss m1_649_17714# vss nfet$197
Xnfet$206_14 m1_15188_21786# m1_15188_21786# vss vss m1_14026_21586# vss nfet$206
Xpfet$182_104 vdd vdd m1_14127_16080# m1_n7513_20152# pfet$182
Xnfet$197_1 m1_9015_17714# vss m1_6116_17343# vss nfet$197
Xpfet$189_2 vdd vdd m1_n1271_25858# m1_n10452_25858# pfet$189
Xpfet$185_13 vdd vdd m1_15188_21786# m1_14556_21786# pfet$185
Xpfet$182_9 vdd vdd m1_8172_15778# m1_5302_17714# pfet$182
Xnfet$217_2 m1_n6788_16080# m1_n6788_16080# m1_n7247_17714# m1_n7247_17714# m1_n6690_16398#
+ vss nfet$217
Xpfet$194_0 vdd vdd m1_n1263_21786# pd1 pfet$194
Xpfet$209_3 vdd vdd vdd m1_n8047_22344# m1_n8283_19850# m1_n8283_19850# pfet$209
Xnfet$194_19 m1_7456_23922# vss m1_8076_24224# vss nfet$194
Xpfet$182_69 vdd vdd m1_20721_15778# m1_17851_17714# pfet$182
Xpfet$182_14 vdd vdd m1_2092_17836# m1_1933_17343# pfet$182
Xpfet$182_25 vdd vdd m1_1709_17518# m1_1119_17714# pfet$182
Xpfet$182_36 vdd vdd m1_6116_17343# m1_9015_17714# pfet$182
Xpfet$182_47 vdd m1_11738_16080# m1_11271_18030# m1_10299_17343# pfet$182
Xpfet$182_58 vdd vdd m1_n3534_17714# m1_n3064_17714# pfet$182
Xnfet$222_0 m1_n9952_24224# m1_n9952_24224# m1_n10308_24542# m1_n10308_24542# m1_n9854_24542#
+ vss nfet$222
Xpfet$207_0 vdd vdd m1_n10796_25662# m1_n10933_25858# pfet$207
Xpfet$200_7 vdd m1_27292_16202# m1_26807_17518# m1_27190_17836# pfet$200
Xnfet$201_5 m1_n7247_17714# vss m1_n6657_17518# vss nfet$201
Xnfet$214_14 m1_22205_20152# m1_22205_20152# m1_n2543_20130# m1_n2543_20130# m1_21039_20470#
+ vss nfet$214
Xnfet$199_5 m1_965_15478# vss m1_8137_20152# vss nfet$199
Xnfet$197_19 m1_n7513_20152# vss m1_1578_16080# vss nfet$197
Xnfet$197_2 m1_6275_17836# m1_7555_16080# m1_7088_18030# vss nfet$197
Xpfet$185_14 vdd vdd m1_19969_21590# m1_19839_21786# pfet$185
Xnfet$206_15 m1_14556_21786# m1_14556_21786# vss vss m1_13394_21586# vss nfet$206
Xpfet$182_105 vdd vdd m1_14258_17518# m1_13668_17714# pfet$182
Xpfet$189_3 vdd vdd m1_1607_24542# m1_n789_25858# pfet$189
Xnfet$217_3 m1_n6172_16202# m1_n6172_16202# vss vss m1_n6690_16398# vss nfet$217
Xpfet$194_1 vdd vdd m1_2254_21786# pd2 pfet$194
Xpfet$187_0 vdd vdd m1_2384_19550# m1_n3534_17714# pfet$187
Xnfet$215_0 m1_35837_22102# vss m1_n7513_20152# vss nfet$215
Xnfet$222_1 m1_n9336_24346# m1_n9336_24346# m1_n8625_26174# m1_n8625_26174# m1_n8389_25502#
+ vss nfet$222
Xpfet$182_15 vdd vdd m1_5302_17714# m1_5761_16080# pfet$182
Xpfet$182_26 vdd vdd m1_4832_17714# m1_5302_17714# pfet$182
Xpfet$182_37 vdd m1_7555_16080# m1_7088_18030# m1_6116_17343# pfet$182
Xpfet$182_48 vdd vdd m1_n3064_17714# m1_n2605_16080# pfet$182
Xpfet$182_59 vdd vdd m1_n2605_16080# m1_n7513_20152# pfet$182
Xpfet$207_1 vdd vdd m1_n10309_25662# m1_n10452_25858# pfet$207
Xnfet$201_6 m1_n7247_17714# vss m1_n7383_17599# vss nfet$201
Xnfet$214_15 m1_17697_15478# m1_17697_15478# m1_n2543_20130# m1_n2543_20130# m1_20407_20470#
+ vss nfet$214
Xnfet$199_6 m1_9015_17714# vss m1_12935_19550# vss nfet$199
Xnfet$197_3 m1_n7513_20152# vss m1_9944_16080# vss nfet$197
Xpfet$185_15 vdd vdd m1_27003_21590# m1_26873_21786# pfet$185
Xnfet$206_16 m1_28624_21786# m1_28624_21786# vss vss m1_27462_21586# vss nfet$206
Xpfet$182_106 vdd vdd m1_14482_17343# m1_17381_17714# pfet$182
Xpfet$189_4 vdd vdd m1_488_21786# m1_n789_25858# pfet$189
Xnfet$217_4 m1_28113_15778# m1_28113_15778# m1_28003_18030# m1_28003_18030# m1_28239_17358#
+ vss nfet$217
Xpfet$194_2 vdd vdd m1_26873_21786# pd9 pfet$194
Xnfet$195_0 m1_n1133_21590# m1_n1133_21590# m1_354_22513# m1_354_22513# m1_n674_21586#
+ vss nfet$195
Xpfet$187_1 vdd vdd m1_4620_20152# m1_n3218_15478# pfet$187
Xnfet$208_0 m1_34843_21786# m1_34843_21786# m1_34093_22102# m1_34093_22102# m1_34329_21430#
+ vss nfet$208
Xnfet$222_2 m1_n8848_25658# m1_n8848_25658# vss vss m1_n8389_25502# vss nfet$222
Xpfet$182_16 vdd vdd m1_3989_15778# m1_1119_17714# pfet$182
Xpfet$182_27 vdd m1_2194_16202# m1_1709_17518# m1_2092_17836# pfet$182
Xpfet$182_38 vdd vdd m1_7088_18030# m1_7198_15778# pfet$182
Xpfet$182_49 vdd m1_n194_15778# m1_n811_16080# m1_n2091_17836# pfet$182
Xpfet$207_2 vdd vdd m1_n9952_24224# m1_n10572_23922# pfet$207
Xnfet$201_7 m1_26217_17714# vss m1_26807_17518# vss nfet$201
Xnfet$214_16 m1_25722_20152# m1_25722_20152# m1_n3206_20274# m1_n3206_20274# m1_24556_20470#
+ vss nfet$214
Xpfet$212_0 vdd vdd vdd m1_n5019_19550# m1_n4485_20152# m1_n4485_20152# pfet$212
Xnfet$199_7 m1_5148_15478# vss m1_11654_20152# vss nfet$199
Xnfet$197_4 m1_10299_17343# m1_10560_16202# m1_10075_17518# vss nfet$197
Xpfet$185_16 vdd vdd m1_29256_21786# m1_28624_21786# pfet$185
Xnfet$206_17 m1_29256_21786# m1_29256_21786# vss vss m1_28094_21586# vss nfet$206
Xpfet$182_107 vdd m1_15921_16080# m1_15454_18030# m1_14482_17343# pfet$182
Xpfet$189_5 vdd vdd m1_326_24346# m1_n7513_20152# pfet$189
Xnfet$217_5 m1_26676_16080# m1_26676_16080# vss vss m1_28239_17358# vss nfet$217
Xnfet$195_1 m1_n1263_21786# m1_n1263_21786# m1_354_22513# m1_354_22513# m1_n42_21586#
+ vss nfet$195
Xpfet$187_2 vdd vdd m1_1103_20152# m1_n7401_15478# pfet$187
Xnfet$208_1 m1_28490_22513# m1_28490_22513# vss vss m1_34329_21430# vss nfet$208
Xnfet$222_3 m1_n9336_24346# m1_n9336_24346# vss vss m1_n9854_24542# vss nfet$222
Xpfet$192_0 vdd m1_31535_19792# vdd m1_17939_22513# pfet$192
Xpfet$182_17 vdd vdd m1_n2091_17836# m1_n2250_17343# pfet$182
Xpfet$182_28 vdd m1_2905_18030# vdd m1_1578_16080# pfet$182
Xpfet$182_39 vdd m1_7088_18030# vdd m1_5761_16080# pfet$182
Xpfet$207_3 vdd vdd m1_n4978_24224# vss pfet$207
Xnfet$201_8 m1_n7513_20152# vss m1_26676_16080# vss nfet$201
Xnfet$195_10 m1_19839_21786# m1_19839_21786# m1_21456_22513# m1_21456_22513# m1_21060_21586#
+ vss nfet$195
Xnfet$214_17 m1_21880_15478# m1_21880_15478# m1_n3206_20274# m1_n3206_20274# m1_23924_20470#
+ vss nfet$214
Xnfet$220_0 m1_n3822_20130# m1_n3822_20130# m1_n4485_20152# m1_n4485_20152# m1_n3724_20470#
+ vss nfet$220
Xpfet$205_0 vdd vdd m1_n8625_26174# m1_n9336_24346# pfet$205
Xnfet$199_8 m1_n7383_17599# vss m1_n1133_19550# vss nfet$199
.ends

.subckt nfet$186 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$176 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$174 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$187 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt nfet$185 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$175 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$173 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$188 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_drive_buffer vss in vdd out
Xnfet$186_0 out out vss m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# m1_4274_n1060#
+ m1_4274_n1060# out m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# vss vss
+ nfet$186
Xpfet$176_0 vdd vdd m1_3466_n454# in pfet$176
Xpfet$174_0 m1_4274_n1060# vdd vdd m1_4274_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ vdd m1_4002_n1060# m1_4002_n1060# pfet$174
Xnfet$187_0 m1_3466_n454# vss m1_4002_n1060# vss nfet$187
Xnfet$185_0 m1_4274_n1060# vss m1_4002_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ m1_4274_n1060# vss m1_4002_n1060# vss nfet$185
Xpfet$175_0 vdd vdd m1_4002_n1060# m1_3466_n454# pfet$175
Xpfet$173_0 out out m1_4274_n1060# vdd m1_4274_n1060# out vdd vdd m1_4274_n1060# out
+ m1_4274_n1060# m1_4274_n1060# out m1_4274_n1060# vdd m1_4274_n1060# vdd m1_4274_n1060#
+ pfet$173
Xnfet$188_0 in vss m1_3466_n454# vss nfet$188
.ends

.subckt pfet$33 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$39 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$34 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$40 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt xp_3_1_MUX$1 S0 S1 VDD VSS OUT_1 C_1 B_1 A_1
Xpfet$33_0 VDD A_1 m1_239_n318# m1_n432_458# pfet$33
Xpfet$33_1 VDD C_1 OUT_1 S1 pfet$33
Xpfet$33_2 VDD B_1 m1_239_n318# S0 pfet$33
Xpfet$33_3 VDD m1_239_n318# OUT_1 m1_n432_n1290# pfet$33
Xnfet$39_0 m1_n432_n1290# C_1 OUT_1 VSS nfet$39
Xnfet$39_1 m1_n432_458# B_1 m1_239_n318# VSS nfet$39
Xnfet$39_2 S1 m1_239_n318# OUT_1 VSS nfet$39
Xnfet$39_3 S0 A_1 m1_239_n318# VSS nfet$39
Xpfet$34_0 VDD VDD m1_n432_n1290# S1 pfet$34
Xpfet$34_1 VDD VDD m1_n432_458# S0 pfet$34
Xnfet$40_0 S1 VSS m1_n432_n1290# VSS nfet$40
Xnfet$40_1 S0 VSS m1_n432_458# VSS nfet$40
.ends

.subckt pfet$217 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$215 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$5 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$3 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$1 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$218 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$216 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$214 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$4 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$2 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt asc_hysteresis_buffer vss in vdd out
Xpfet$217_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$217
Xpfet$215_0 vdd vdd m1_884_42# m1_348_648# pfet$215
Xnfet$5_0 m1_1156_42# vss m1_884_42# vss nfet$5
Xnfet$3_0 in vss m1_348_648# vss nfet$3
Xnfet$1_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$1
Xpfet$218_0 vdd vdd m1_884_42# m1_1156_42# pfet$218
Xpfet$216_0 vdd vdd m1_348_648# in pfet$216
Xpfet$214_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd
+ m1_884_42# m1_884_42# pfet$214
Xnfet$4_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$4
Xnfet$2_0 m1_348_648# vss m1_884_42# vss nfet$2
.ends

.subckt nfet$15 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$1 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$17 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$8 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$6 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$9 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$14 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$20 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$13 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$4 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$7 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$12 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$11 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$2 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$10 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$5 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$18 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$9 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$16 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$7 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$15 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$14 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$8 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$13 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$12 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$3 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$6 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$11 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$10 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt nfet$19 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_lock_detector_20250826 ref vdd div lock vss
Xnfet$15_10 m1_12790_7868# vss m1_15618_7156# vss nfet$15
Xpfet$1_6 vdd vdd m1_2446_5099# m1_208_7868# pfet$1
Xnfet$17_0 div m1_n4030_5270# vss vss nfet$17
Xnfet$15_11 m1_15979_5220# vss m1_16599_5522# vss nfet$15
Xpfet$1_7 vdd vdd m1_2446_1478# m1_208_n340# pfet$1
Xpfet$8_0 m1_n10260_7868# m1_n10260_7868# m1_n11408_4493# vdd m1_n11408_4493# m1_n10260_7868#
+ vdd vdd m1_n11408_4493# m1_n10260_7868# m1_n11408_4493# m1_n11408_4493# m1_n10260_7868#
+ m1_n11408_4493# vdd m1_n11408_4493# vdd m1_n11408_4493# pfet$8
Xnfet$17_1 m1_n6066_7868# vss m1_n4030_5270# vss nfet$17
Xnfet$15_12 m1_15618_7156# vss m1_15755_6960# vss nfet$15
Xpfet$8_1 m1_n6066_7868# m1_n6066_7868# m1_n7214_4493# vdd m1_n7214_4493# m1_n6066_7868#
+ vdd vdd m1_n7214_4493# m1_n6066_7868# m1_n7214_4493# m1_n7214_4493# m1_n6066_7868#
+ m1_n7214_4493# vdd m1_n7214_4493# vdd m1_n7214_4493# pfet$8
Xnfet$15_13 ref vss m1_16242_6960# vss nfet$15
Xpfet$8_2 m1_n14454_7868# m1_n14454_7868# m1_n15602_4493# vdd m1_n15602_4493# m1_n14454_7868#
+ vdd vdd m1_n15602_4493# m1_n14454_7868# m1_n15602_4493# m1_n15602_4493# m1_n14454_7868#
+ m1_n15602_4493# vdd m1_n15602_4493# vdd m1_n15602_4493# pfet$8
Xnfet$15_0 m1_15979_2344# vss m1_16599_2028# vss nfet$15
Xpfet$6_0 vdd m1_16599_2028# m1_17703_788# m1_15618_394# pfet$6
Xnfet$9_0 m1_n6066_7868# m1_n6066_7868# vss m1_n7214_4493# m1_n7214_4493# m1_n6066_7868#
+ vss m1_n7214_4493# m1_n7214_4493# m1_n7214_4493# m1_n6066_7868# m1_n7214_4493# m1_n7214_4493#
+ m1_n6066_7868# vss m1_n7214_4493# vss vss nfet$9
Xnfet$15_1 m1_15618_394# vss m1_15755_n208# vss nfet$15
Xpfet$14_0 vdd m1_19675_2344# vdd m1_19469_1832# pfet$14
Xpfet$6_1 vdd m1_16242_n208# m1_15979_2344# m1_15755_n208# pfet$6
Xnfet$9_1 m1_n14454_7868# m1_n14454_7868# vss m1_n15602_4493# m1_n15602_4493# m1_n14454_7868#
+ vss m1_n15602_4493# m1_n15602_4493# m1_n15602_4493# m1_n14454_7868# m1_n15602_4493#
+ m1_n15602_4493# m1_n14454_7868# vss m1_n15602_4493# vss vss nfet$9
Xnfet$15_2 m1_n2336_5099# vss m1_16242_n208# vss nfet$15
Xpfet$14_1 vdd vdd m1_19675_2344# m1_19469_4920# pfet$14
Xnfet$20_0 m1_19675_2344# vss lock vss nfet$20
Xpfet$6_2 vdd m1_15979_2344# m1_16243_1828# m1_15618_394# pfet$6
Xnfet$9_2 m1_n10260_7868# m1_n10260_7868# vss m1_n11408_4493# m1_n11408_4493# m1_n10260_7868#
+ vss m1_n11408_4493# m1_n11408_4493# m1_n11408_4493# m1_n10260_7868# m1_n11408_4493#
+ m1_n11408_4493# m1_n10260_7868# vss m1_n11408_4493# vss vss nfet$9
Xnfet$15_3 m1_17926_34# vss m1_18496_1828# vss nfet$15
Xnfet$13_0 m1_15755_n208# m1_16599_2028# m1_17703_788# vss nfet$13
Xpfet$6_3 vdd m1_17703_788# m1_18496_1828# m1_15755_n208# pfet$6
Xpfet$4_0 m1_7448_n340# vdd vdd m1_7448_n340# m1_7176_n340# m1_7176_n340# m1_7448_n340#
+ vdd m1_7176_n340# m1_7176_n340# pfet$4
Xnfet$15_4 m1_12790_n340# vss m1_15618_394# vss nfet$15
Xnfet$13_1 m1_15618_394# m1_16242_n208# m1_15979_2344# vss nfet$13
Xnfet$7_0 m1_10834_1478# vss m1_11370_n340# vss nfet$7
Xpfet$6_4 vdd m1_17703_6956# m1_18496_5840# m1_15755_6960# pfet$6
Xpfet$12_0 vdd vdd vdd m1_n3798_6028# div div pfet$12
Xpfet$4_1 m1_11642_n340# vdd vdd m1_11642_n340# m1_11370_n340# m1_11370_n340# m1_11642_n340#
+ vdd m1_11370_n340# m1_11370_n340# pfet$4
Xnfet$7_1 m1_2446_1478# vss m1_2982_n340# vss nfet$7
Xnfet$15_5 vss vss m1_17215_2028# vss nfet$15
Xnfet$13_2 m1_15618_394# m1_17703_788# m1_18496_1828# vss nfet$13
Xpfet$12_1 vdd m1_n4030_5270# m1_n4030_5270# m1_n3798_6028# m1_n6066_7868# m1_n6066_7868#
+ pfet$12
Xpfet$6_5 vdd m1_15979_5220# m1_16243_5840# m1_15618_7156# pfet$6
Xpfet$4_2 m1_3254_n340# vdd vdd m1_3254_n340# m1_2982_n340# m1_2982_n340# m1_3254_n340#
+ vdd m1_2982_n340# m1_2982_n340# pfet$4
Xnfet$7_2 m1_6640_1478# vss m1_7176_n340# vss nfet$7
Xnfet$13_3 m1_15755_n208# m1_15979_2344# m1_16243_1828# vss nfet$13
Xnfet$15_6 m1_17926_34# vss m1_19469_1832# vss nfet$15
Xnfet$11_0 m1_n7214_4493# vss m1_n7486_4493# m1_n7486_4493# m1_n7486_4493# m1_n7214_4493#
+ m1_n7214_4493# vss m1_n7486_4493# vss nfet$11
Xpfet$6_6 vdd m1_16599_5522# m1_17703_6956# m1_15618_7156# pfet$6
Xpfet$4_3 m1_n940_n340# vdd vdd m1_n940_n340# m1_n1212_n340# m1_n1212_n340# m1_n940_n340#
+ vdd m1_n1212_n340# m1_n1212_n340# pfet$4
Xpfet$2_0 vdd vdd m1_7176_n340# m1_6640_1478# pfet$2
Xnfet$7_3 m1_n1748_1478# vss m1_n1212_n340# vss nfet$7
Xnfet$15_7 vss vss m1_17215_5644# vss nfet$15
Xnfet$11_1 m1_n15602_4493# vss m1_n15874_4493# m1_n15874_4493# m1_n15874_4493# m1_n15602_4493#
+ m1_n15602_4493# vss m1_n15874_4493# vss nfet$11
Xnfet$13_4 m1_15618_7156# m1_17703_6956# m1_18496_5840# vss nfet$13
Xpfet$6_7 vdd m1_16242_6960# m1_15979_5220# m1_15755_6960# pfet$6
Xpfet$10_0 vdd vdd m1_n11680_4493# m1_n12216_5099# pfet$10
Xpfet$2_1 vdd vdd m1_11370_n340# m1_10834_1478# pfet$2
Xpfet$4_4 m1_n940_4493# vdd vdd m1_n940_4493# m1_n1212_4493# m1_n1212_4493# m1_n940_4493#
+ vdd m1_n1212_4493# m1_n1212_4493# pfet$4
Xnfet$7_4 m1_10834_5099# vss m1_11370_4493# vss nfet$7
Xnfet$13_5 m1_15755_6960# m1_15979_5220# m1_16243_5840# vss nfet$13
Xnfet$15_8 m1_17926_7472# vss m1_19469_4920# vss nfet$15
Xnfet$11_2 m1_n11408_4493# vss m1_n11680_4493# m1_n11680_4493# m1_n11680_4493# m1_n11408_4493#
+ m1_n11408_4493# vss m1_n11680_4493# vss nfet$11
Xpfet$4_5 m1_11642_4493# vdd vdd m1_11642_4493# m1_11370_4493# m1_11370_4493# m1_11642_4493#
+ vdd m1_11370_4493# m1_11370_4493# pfet$4
Xpfet$10_1 vdd vdd m1_n7486_4493# m1_n8022_5099# pfet$10
Xnfet$15_9 m1_17926_7472# vss m1_18496_5840# vss nfet$15
Xpfet$2_2 vdd vdd m1_2982_n340# m1_2446_1478# pfet$2
Xnfet$7_5 m1_6640_5099# vss m1_7176_4493# vss nfet$7
Xnfet$13_6 m1_15618_7156# m1_16242_6960# m1_15979_5220# vss nfet$13
Xpfet$5_10 vdd vdd m1_15618_7156# m1_12790_7868# pfet$5
Xpfet$10_2 vdd vdd m1_n15874_4493# m1_n16410_5099# pfet$10
Xpfet$4_6 m1_3254_4493# vdd vdd m1_3254_4493# m1_2982_4493# m1_2982_4493# m1_3254_4493#
+ vdd m1_2982_4493# m1_2982_4493# pfet$4
Xpfet$2_3 vdd vdd m1_n1212_n340# m1_n1748_1478# pfet$2
Xnfet$7_6 m1_n1748_5099# vss m1_n1212_4493# vss nfet$7
Xnfet$13_7 m1_15755_6960# m1_16599_5522# m1_17703_6956# vss nfet$13
Xpfet$4_7 m1_7448_4493# vdd vdd m1_7448_4493# m1_7176_4493# m1_7176_4493# m1_7448_4493#
+ vdd m1_7176_4493# m1_7176_4493# pfet$4
Xpfet$5_11 vdd vdd m1_16599_5522# m1_15979_5220# pfet$5
Xpfet$2_4 vdd vdd m1_n1212_4493# m1_n1748_5099# pfet$2
Xnfet$7_7 m1_2446_5099# vss m1_2982_4493# vss nfet$7
Xpfet$5_12 vdd vdd m1_16242_6960# ref pfet$5
Xpfet$2_5 vdd vdd m1_2982_4493# m1_2446_5099# pfet$2
Xpfet$5_13 vdd vdd m1_15755_6960# m1_15618_7156# pfet$5
Xpfet$2_6 vdd vdd m1_7176_4493# m1_6640_5099# pfet$2
Xnfet$18_0 m1_n4030_5270# vss m1_n2336_5099# vss nfet$18
Xpfet$9_0 m1_n11408_4493# vdd vdd m1_n11408_4493# m1_n11680_4493# m1_n11680_4493#
+ m1_n11408_4493# vdd m1_n11680_4493# m1_n11680_4493# pfet$9
Xpfet$2_7 vdd vdd m1_11370_4493# m1_10834_5099# pfet$2
Xpfet$9_1 m1_n7214_4493# vdd vdd m1_n7214_4493# m1_n7486_4493# m1_n7486_4493# m1_n7214_4493#
+ vdd m1_n7486_4493# m1_n7486_4493# pfet$9
Xpfet$9_2 m1_n15602_4493# vdd vdd m1_n15602_4493# m1_n15874_4493# m1_n15874_4493#
+ m1_n15602_4493# vdd m1_n15874_4493# m1_n15874_4493# pfet$9
Xnfet$16_0 m1_n14454_7868# vss m1_n12216_5099# vss nfet$16
Xpfet$7_0 vdd m1_17926_34# vdd m1_17703_788# pfet$7
Xnfet$16_1 div vss m1_n16410_5099# vss nfet$16
Xpfet$15_0 vdd vdd lock m1_19675_2344# pfet$15
Xpfet$7_1 vdd vdd m1_17926_34# m1_17215_2028# pfet$7
Xnfet$16_2 m1_n10260_7868# vss m1_n8022_5099# vss nfet$16
Xpfet$7_2 vdd m1_16243_1828# vdd m1_17215_2028# pfet$7
Xnfet$14_0 m1_17215_2028# m1_17215_2028# m1_17926_34# m1_17926_34# m1_18162_712# vss
+ nfet$14
Xpfet$7_3 vdd vdd m1_16243_1828# m1_16599_2028# pfet$7
Xpfet$5_0 vdd vdd m1_16599_2028# m1_15979_2344# pfet$5
Xnfet$14_1 m1_17703_788# m1_17703_788# vss vss m1_18162_712# vss nfet$14
Xnfet$8_0 m1_3254_n340# vss m1_2982_n340# m1_2982_n340# m1_2982_n340# m1_3254_n340#
+ m1_3254_n340# vss m1_2982_n340# vss nfet$8
Xpfet$13_0 vdd vdd m1_n2336_5099# m1_n4030_5270# pfet$13
Xpfet$5_1 vdd vdd m1_16242_n208# m1_n2336_5099# pfet$5
Xpfet$7_4 vdd m1_16243_5840# vdd m1_17215_5644# pfet$7
Xnfet$8_1 m1_7448_n340# vss m1_7176_n340# m1_7176_n340# m1_7176_n340# m1_7448_n340#
+ m1_7448_n340# vss m1_7176_n340# vss nfet$8
Xnfet$14_2 m1_16599_2028# m1_16599_2028# m1_16243_1828# m1_16243_1828# m1_16697_1672#
+ vss nfet$14
Xpfet$7_5 vdd vdd m1_16243_5840# m1_16599_5522# pfet$7
Xpfet$5_2 vdd vdd m1_15755_n208# m1_15618_394# pfet$5
Xnfet$8_2 m1_11642_n340# vss m1_11370_n340# m1_11370_n340# m1_11370_n340# m1_11642_n340#
+ m1_11642_n340# vss m1_11370_n340# vss nfet$8
Xnfet$12_0 m1_8596_n340# vss m1_10834_1478# vss nfet$12
Xnfet$14_3 m1_17215_2028# m1_17215_2028# vss vss m1_16697_1672# vss nfet$14
Xpfet$7_6 vdd m1_17926_7472# vdd m1_17703_6956# pfet$7
Xpfet$5_3 vdd vdd m1_18496_1828# m1_17926_34# pfet$5
Xpfet$3_0 m1_8596_n340# m1_8596_n340# m1_7448_n340# vdd m1_7448_n340# m1_8596_n340#
+ vdd vdd m1_7448_n340# m1_8596_n340# m1_7448_n340# m1_7448_n340# m1_8596_n340# m1_7448_n340#
+ vdd m1_7448_n340# vdd m1_7448_n340# pfet$3
Xnfet$6_0 m1_8596_n340# m1_8596_n340# vss m1_7448_n340# m1_7448_n340# m1_8596_n340#
+ vss m1_7448_n340# m1_7448_n340# m1_7448_n340# m1_8596_n340# m1_7448_n340# m1_7448_n340#
+ m1_8596_n340# vss m1_7448_n340# vss vss nfet$6
Xnfet$8_3 m1_n940_n340# vss m1_n1212_n340# m1_n1212_n340# m1_n1212_n340# m1_n940_n340#
+ m1_n940_n340# vss m1_n1212_n340# vss nfet$8
Xnfet$14_4 m1_17215_5644# m1_17215_5644# vss vss m1_16697_5840# vss nfet$14
Xpfet$7_7 vdd vdd m1_17926_7472# m1_17215_5644# pfet$7
Xnfet$12_1 m1_4402_n340# vss m1_6640_1478# vss nfet$12
Xpfet$11_0 vdd vdd m1_n8022_5099# m1_n10260_7868# pfet$11
Xpfet$5_4 vdd vdd m1_15618_394# m1_12790_n340# pfet$5
Xnfet$8_4 m1_11642_4493# vss m1_11370_4493# m1_11370_4493# m1_11370_4493# m1_11642_4493#
+ m1_11642_4493# vss m1_11370_4493# vss nfet$8
Xpfet$3_1 m1_12790_n340# m1_12790_n340# m1_11642_n340# vdd m1_11642_n340# m1_12790_n340#
+ vdd vdd m1_11642_n340# m1_12790_n340# m1_11642_n340# m1_11642_n340# m1_12790_n340#
+ m1_11642_n340# vdd m1_11642_n340# vdd m1_11642_n340# pfet$3
Xnfet$14_5 m1_16599_5522# m1_16599_5522# m1_16243_5840# m1_16243_5840# m1_16697_5840#
+ vss nfet$14
Xnfet$6_1 m1_4402_n340# m1_4402_n340# vss m1_3254_n340# m1_3254_n340# m1_4402_n340#
+ vss m1_3254_n340# m1_3254_n340# m1_3254_n340# m1_4402_n340# m1_3254_n340# m1_3254_n340#
+ m1_4402_n340# vss m1_3254_n340# vss vss nfet$6
Xnfet$12_2 ref vss m1_n1748_1478# vss nfet$12
Xpfet$11_1 vdd vdd m1_n16410_5099# div pfet$11
Xpfet$5_5 vdd vdd m1_17215_2028# vss pfet$5
Xpfet$3_2 m1_4402_n340# m1_4402_n340# m1_3254_n340# vdd m1_3254_n340# m1_4402_n340#
+ vdd vdd m1_3254_n340# m1_4402_n340# m1_3254_n340# m1_3254_n340# m1_4402_n340# m1_3254_n340#
+ vdd m1_3254_n340# vdd m1_3254_n340# pfet$3
Xnfet$8_5 m1_7448_4493# vss m1_7176_4493# m1_7176_4493# m1_7176_4493# m1_7448_4493#
+ m1_7448_4493# vss m1_7176_4493# vss nfet$8
Xnfet$14_6 m1_17215_5644# m1_17215_5644# m1_17926_7472# m1_17926_7472# m1_18162_6800#
+ vss nfet$14
Xnfet$6_2 m1_12790_n340# m1_12790_n340# vss m1_11642_n340# m1_11642_n340# m1_12790_n340#
+ vss m1_11642_n340# m1_11642_n340# m1_11642_n340# m1_12790_n340# m1_11642_n340# m1_11642_n340#
+ m1_12790_n340# vss m1_11642_n340# vss vss nfet$6
Xnfet$12_3 m1_n2336_5099# vss m1_n1748_5099# vss nfet$12
Xpfet$11_2 vdd vdd m1_n12216_5099# m1_n14454_7868# pfet$11
Xnfet$10_0 m1_n8022_5099# vss m1_n7486_4493# vss nfet$10
Xpfet$5_6 vdd vdd m1_19469_1832# m1_17926_34# pfet$5
Xnfet$8_6 m1_n940_4493# vss m1_n1212_4493# m1_n1212_4493# m1_n1212_4493# m1_n940_4493#
+ m1_n940_4493# vss m1_n1212_4493# vss nfet$8
Xpfet$1_0 vdd vdd m1_6640_1478# m1_4402_n340# pfet$1
Xpfet$3_3 m1_208_n340# m1_208_n340# m1_n940_n340# vdd m1_n940_n340# m1_208_n340# vdd
+ vdd m1_n940_n340# m1_208_n340# m1_n940_n340# m1_n940_n340# m1_208_n340# m1_n940_n340#
+ vdd m1_n940_n340# vdd m1_n940_n340# pfet$3
Xnfet$14_7 m1_17703_6956# m1_17703_6956# vss vss m1_18162_6800# vss nfet$14
Xnfet$12_4 m1_8596_7868# vss m1_10834_5099# vss nfet$12
Xnfet$6_3 m1_208_n340# m1_208_n340# vss m1_n940_n340# m1_n940_n340# m1_208_n340# vss
+ m1_n940_n340# m1_n940_n340# m1_n940_n340# m1_208_n340# m1_n940_n340# m1_n940_n340#
+ m1_208_n340# vss m1_n940_n340# vss vss nfet$6
Xnfet$10_1 m1_n16410_5099# vss m1_n15874_4493# vss nfet$10
Xpfet$3_4 m1_208_7868# m1_208_7868# m1_n940_4493# vdd m1_n940_4493# m1_208_7868# vdd
+ vdd m1_n940_4493# m1_208_7868# m1_n940_4493# m1_n940_4493# m1_208_7868# m1_n940_4493#
+ vdd m1_n940_4493# vdd m1_n940_4493# pfet$3
Xpfet$5_7 vdd vdd m1_17215_5644# vss pfet$5
Xnfet$8_7 m1_3254_4493# vss m1_2982_4493# m1_2982_4493# m1_2982_4493# m1_3254_4493#
+ m1_3254_4493# vss m1_2982_4493# vss nfet$8
Xpfet$1_1 vdd vdd m1_10834_1478# m1_8596_n340# pfet$1
Xnfet$6_4 m1_12790_7868# m1_12790_7868# vss m1_11642_4493# m1_11642_4493# m1_12790_7868#
+ vss m1_11642_4493# m1_11642_4493# m1_11642_4493# m1_12790_7868# m1_11642_4493# m1_11642_4493#
+ m1_12790_7868# vss m1_11642_4493# vss vss nfet$6
Xnfet$12_5 m1_4402_7868# vss m1_6640_5099# vss nfet$12
Xnfet$10_2 m1_n12216_5099# vss m1_n11680_4493# vss nfet$10
Xpfet$5_8 vdd vdd m1_19469_4920# m1_17926_7472# pfet$5
Xpfet$3_5 m1_12790_7868# m1_12790_7868# m1_11642_4493# vdd m1_11642_4493# m1_12790_7868#
+ vdd vdd m1_11642_4493# m1_12790_7868# m1_11642_4493# m1_11642_4493# m1_12790_7868#
+ m1_11642_4493# vdd m1_11642_4493# vdd m1_11642_4493# pfet$3
Xnfet$6_5 m1_8596_7868# m1_8596_7868# vss m1_7448_4493# m1_7448_4493# m1_8596_7868#
+ vss m1_7448_4493# m1_7448_4493# m1_7448_4493# m1_8596_7868# m1_7448_4493# m1_7448_4493#
+ m1_8596_7868# vss m1_7448_4493# vss vss nfet$6
Xpfet$1_2 vdd vdd m1_n1748_1478# ref pfet$1
Xnfet$12_6 m1_208_n340# vss m1_2446_1478# vss nfet$12
Xpfet$3_6 m1_4402_7868# m1_4402_7868# m1_3254_4493# vdd m1_3254_4493# m1_4402_7868#
+ vdd vdd m1_3254_4493# m1_4402_7868# m1_3254_4493# m1_3254_4493# m1_4402_7868# m1_3254_4493#
+ vdd m1_3254_4493# vdd m1_3254_4493# pfet$3
Xpfet$5_9 vdd vdd m1_18496_5840# m1_17926_7472# pfet$5
Xpfet$1_3 vdd vdd m1_n1748_5099# m1_n2336_5099# pfet$1
Xnfet$6_6 m1_208_7868# m1_208_7868# vss m1_n940_4493# m1_n940_4493# m1_208_7868# vss
+ m1_n940_4493# m1_n940_4493# m1_n940_4493# m1_208_7868# m1_n940_4493# m1_n940_4493#
+ m1_208_7868# vss m1_n940_4493# vss vss nfet$6
Xnfet$12_7 m1_208_7868# vss m1_2446_5099# vss nfet$12
Xnfet$19_0 m1_19469_4920# m1_19469_4920# m1_19675_2344# m1_19675_2344# m1_19911_1672#
+ vss nfet$19
Xpfet$3_7 m1_8596_7868# m1_8596_7868# m1_7448_4493# vdd m1_7448_4493# m1_8596_7868#
+ vdd vdd m1_7448_4493# m1_8596_7868# m1_7448_4493# m1_7448_4493# m1_8596_7868# m1_7448_4493#
+ vdd m1_7448_4493# vdd m1_7448_4493# pfet$3
Xnfet$6_7 m1_4402_7868# m1_4402_7868# vss m1_3254_4493# m1_3254_4493# m1_4402_7868#
+ vss m1_3254_4493# m1_3254_4493# m1_3254_4493# m1_4402_7868# m1_3254_4493# m1_3254_4493#
+ m1_4402_7868# vss m1_3254_4493# vss vss nfet$6
Xpfet$1_4 vdd vdd m1_6640_5099# m1_4402_7868# pfet$1
Xnfet$19_1 m1_19469_1832# m1_19469_1832# vss vss m1_19911_1672# vss nfet$19
Xpfet$1_5 vdd vdd m1_10834_5099# m1_8596_7868# pfet$1
.ends

.subckt asc_dual_psd_def_20250809$1 vdd vss pd1 pd2 pd3 pd4 pd5 pd6 pd7 pd8 pd9 fout
+ sd1 sd2 sd3 sd4 sd5 sd6 sd7 sd8 sd9 fin define
Xpfet$185_17 vdd vdd m1_25739_21786# m1_25107_21786# pfet$185
Xpfet$182_108 vdd vdd m1_15454_18030# m1_15564_15778# pfet$182
Xpfet$189_6 vdd vdd m1_n290_24224# m1_n910_23922# pfet$189
Xnfet$197_5 m1_10458_17836# m1_11738_16080# m1_11271_18030# vss nfet$197
Xnfet$198_10 m1_21590_21786# vss m1_22222_21786# vss nfet$198
Xnfet$217_6 m1_27292_16202# m1_27292_16202# vss vss m1_26774_16398# vss nfet$217
Xnfet$195_2 m1_9288_21786# m1_9288_21786# m1_9645_21447# m1_9645_21447# m1_10509_21586#
+ vss nfet$195
Xpfet$187_3 vdd vdd m1_5901_19550# m1_649_17714# pfet$187
Xnfet$222_4 m1_n4978_24224# m1_n4978_24224# m1_n10452_25858# m1_n10452_25858# m1_n4880_24542#
+ vss nfet$222
Xnfet$208_2 m1_9645_21447# m1_9645_21447# vss vss m1_30492_21430# vss nfet$208
Xpfet$182_18 vdd m1_1119_17714# vdd m1_2194_16202# pfet$182
Xpfet$182_29 vdd vdd m1_1578_16080# m1_n7513_20152# pfet$182
Xpfet$207_4 vdd vdd m1_n5571_25662# m1_n10452_25858# pfet$207
Xpfet$192_1 vdd vdd m1_30256_19792# m1_21456_22513# pfet$192
Xnfet$201_9 m1_n10452_25858# vss m1_27031_17343# vss nfet$201
Xpfet$185_0 vdd vdd m1_n1133_21590# m1_n1263_21786# pfet$185
Xnfet$195_11 m1_19969_21590# m1_19969_21590# m1_21456_22513# m1_21456_22513# m1_20428_21586#
+ vss nfet$195
Xnfet$213_0 m1_7198_15778# m1_7198_15778# m1_7088_18030# m1_7088_18030# m1_7324_17358#
+ vss nfet$213
Xnfet$220_1 m1_n1927_20274# m1_n1927_20274# vss vss m1_n2445_20470# vss nfet$220
Xpfet$205_1 vdd m1_n8625_26174# vdd m1_n8848_25658# pfet$205
Xnfet$199_9 m1_25747_17714# vss m1_27003_19550# vss nfet$199
Xpfet$182_109 vdd vdd m1_10299_17343# m1_13198_17714# pfet$182
Xpfet$189_7 vdd vdd m1_32330_25662# m1_32193_25858# pfet$189
Xnfet$197_6 m1_6116_17343# vss m1_6275_17836# vss nfet$197
Xnfet$217_7 m1_26676_16080# m1_26676_16080# m1_26217_17714# m1_26217_17714# m1_26774_16398#
+ vss nfet$217
Xnfet$195_3 m1_9418_21590# m1_9418_21590# m1_9645_21447# m1_9645_21447# m1_9877_21586#
+ vss nfet$195
Xnfet$198_11 m1_18073_21786# vss m1_18705_21786# vss nfet$198
Xpfet$187_4 vdd vdd m1_12935_19550# m1_9015_17714# pfet$187
Xnfet$208_3 m1_7388_22513# m1_7388_22513# m1_30256_22102# m1_30256_22102# m1_30492_21430#
+ vss nfet$208
Xpfet$182_19 vdd m1_3015_15778# m1_2194_16202# m1_1933_17343# pfet$182
Xnfet$222_5 m1_n4362_24346# m1_n4362_24346# vss vss m1_n4880_24542# vss nfet$222
Xpfet$207_5 vdd vdd m1_n4847_25662# m1_n10452_25858# pfet$207
Xnfet$193_0 m1_4509_24346# m1_4509_24346# vss vss m1_3991_24542# vss nfet$193
Xpfet$192_2 vdd m1_30256_19792# vdd m1_24973_22513# pfet$192
Xpfet$185_1 vdd vdd m1_11671_21786# m1_11039_21786# pfet$185
Xnfet$195_12 m1_16322_21786# m1_16322_21786# m1_17939_22513# m1_17939_22513# m1_17543_21586#
+ vss nfet$195
Xnfet$213_1 m1_5761_16080# m1_5761_16080# vss vss m1_7324_17358# vss nfet$213
Xnfet$220_2 m1_n3206_20274# m1_n3206_20274# vss vss m1_n3724_20470# vss nfet$220
Xnfet$206_0 m1_11039_21786# m1_11039_21786# vss vss m1_9877_21586# vss nfet$206
Xpfet$205_2 vdd m1_n3651_26174# vdd m1_n4978_24224# pfet$205
Xpfet$210_0 vdd m1_n6380_21786# m1_n6380_21786# m1_n5019_19550# m1_n5227_20152# m1_n5227_20152#
+ pfet$210
Xnfet$197_7 m1_9485_17714# vss m1_10075_17518# vss nfet$197
Xpfet$189_8 vdd vdd m1_33174_24224# m1_32554_23922# pfet$189
Xpfet$181_110 vdd m1_11903_24542# vdd m1_12875_24346# pfet$181
Xnfet$198_12 m1_14556_21786# vss m1_15188_21786# vss nfet$198
Xpfet$187_5 vdd vdd m1_8137_20152# m1_965_15478# pfet$187
Xnfet$195_4 m1_5901_21590# m1_5901_21590# m1_7388_22513# m1_7388_22513# m1_6360_21586#
+ vss nfet$195
Xnfet$222_6 m1_n4978_24224# m1_n4978_24224# vss vss m1_n3415_25502# vss nfet$222
Xnfet$193_1 m1_3893_24224# m1_3893_24224# m1_3537_24542# m1_3537_24542# m1_3991_24542#
+ vss nfet$193
Xpfet$192_3 vdd vdd m1_34843_21786# m1_34093_19792# pfet$192
Xpfet$207_6 vdd vdd m1_n4623_25487# fin pfet$207
Xpfet$185_2 vdd vdd m1_12935_21590# m1_12805_21786# pfet$185
Xnfet$195_13 m1_16452_21590# m1_16452_21590# m1_17939_22513# m1_17939_22513# m1_16911_21586#
+ vss nfet$195
Xnfet$213_2 m1_9944_16080# m1_9944_16080# vss vss m1_11507_17358# vss nfet$213
Xnfet$220_3 m1_n6973_21481# m1_n6973_21481# m1_n6839_20152# m1_n6839_20152# m1_n6282_20470#
+ vss nfet$220
Xpfet$205_3 vdd vdd m1_n3651_26174# m1_n3541_23922# pfet$205
Xnfet$206_1 m1_11671_21786# m1_11671_21786# vss vss m1_10509_21586# vss nfet$206
Xpfet$183_30 vdd vdd vdd m1_17539_22402# m1_16322_21786# m1_16322_21786# pfet$183
Xpfet$190_0 vdd vdd m1_n646_24542# m1_n290_24224# pfet$190
Xpfet$210_1 vdd vdd vdd m1_n5019_22344# m1_n4485_21904# m1_n4485_21904# pfet$210
Xpfet$203_0 vdd m1_n10309_25662# m1_n10572_23922# m1_n10796_25662# pfet$203
Xnfet$201_10 m1_26217_17714# vss m1_29087_15778# vss nfet$201
Xnfet$197_8 m1_7555_16080# vss m1_7198_15778# vss nfet$197
Xpfet$189_9 vdd vdd m1_28624_21786# m1_32675_25947# pfet$189
Xpfet$181_100 vdd vdd m1_29607_24346# m1_n7513_20152# pfet$181
Xnfet$198_13 m1_16322_21786# vss m1_16452_21590# vss nfet$198
Xnfet$229_0 m1_n6839_20152# vss m1_n8145_21908# vss nfet$229
Xnfet$195_5 m1_2254_21786# m1_2254_21786# m1_3871_22513# m1_3871_22513# m1_3475_21586#
+ vss nfet$195
Xpfet$187_6 vdd vdd m1_9418_19550# m1_4832_17714# pfet$187
Xnfet$193_2 m1_4997_25658# m1_4997_25658# vss vss m1_5456_25502# vss nfet$193
Xnfet$222_7 m1_n3541_23922# m1_n3541_23922# m1_n3651_26174# m1_n3651_26174# m1_n3415_25502#
+ vss nfet$222
Xpfet$192_4 vdd m1_34093_19792# vdd m1_32818_20470# pfet$192
Xpfet$207_7 vdd vdd m1_n3541_23922# m1_n3184_24224# pfet$207
Xpfet$185_3 vdd vdd m1_9418_21590# m1_9288_21786# pfet$185
Xnfet$195_14 m1_12805_21786# m1_12805_21786# m1_14422_22513# m1_14422_22513# m1_14026_21586#
+ vss nfet$195
Xnfet$213_3 m1_11381_15778# m1_11381_15778# m1_11271_18030# m1_11271_18030# m1_11507_17358#
+ vss nfet$213
Xnfet$220_4 m1_2590_19404# m1_2590_19404# vss vss m1_n2445_21430# vss nfet$220
Xnfet$206_2 m1_8154_21786# m1_8154_21786# vss vss m1_6992_21586# vss nfet$206
Xpfet$183_31 vdd vdd vdd m1_27462_22102# m1_27003_21590# m1_27003_21590# pfet$183
Xpfet$183_20 vdd vdd vdd m1_20428_22102# m1_19969_21590# m1_19969_21590# pfet$183
Xpfet$190_1 vdd m1_n789_25858# vdd m1_814_25658# pfet$190
Xpfet$183_0 vdd vdd vdd m1_n674_22102# m1_n1133_21590# m1_n1133_21590# pfet$183
Xpfet$205_4 vdd m1_n10452_25858# vdd m1_n4362_24346# pfet$205
Xnfet$211_0 m1_34093_22102# vss fout vss nfet$211
Xpfet$210_2 vdd m1_n5764_21786# m1_n5764_21786# m1_n5019_22344# m1_n5227_21418# m1_n5227_21418#
+ pfet$210
Xpfet$203_1 vdd m1_n9952_24224# m1_n8848_25658# m1_n10933_25858# pfet$203
Xnfet$201_11 m1_27031_17343# vss m1_27190_17836# vss nfet$201
Xnfet$197_9 sd5 vss m1_9331_15478# vss nfet$197
Xpfet$181_101 vdd vdd m1_28010_25858# m1_21590_21786# pfet$181
Xnfet$198_14 m1_19839_21786# vss m1_19969_21590# vss nfet$198
Xnfet$195_6 m1_2384_21590# m1_2384_21590# m1_3871_22513# m1_3871_22513# m1_2843_21586#
+ vss nfet$195
Xpfet$187_7 vdd vdd m1_11654_20152# m1_5148_15478# pfet$187
Xpfet$192_5 vdd vdd m1_34093_19792# m1_32818_21586# pfet$192
Xnfet$193_3 m1_4509_24346# m1_4509_24346# m1_3394_25858# m1_3394_25858# m1_5456_25502#
+ vss nfet$193
Xpfet$207_8 vdd vdd m1_n2567_23922# m1_n7320_25516# pfet$207
Xpfet$185_4 vdd vdd m1_8154_21786# m1_7522_21786# pfet$185
Xnfet$195_15 m1_26873_21786# m1_26873_21786# m1_28490_22513# m1_28490_22513# m1_28094_21586#
+ vss nfet$195
Xnfet$213_4 m1_10560_16202# m1_10560_16202# vss vss m1_10042_16398# vss nfet$213
Xnfet$220_5 m1_6107_19404# m1_6107_19404# m1_n5227_21418# m1_n5227_21418# m1_n2445_21430#
+ vss nfet$220
Xnfet$206_3 m1_7522_21786# m1_7522_21786# vss vss m1_6360_21586# vss nfet$206
Xpfet$183_32 vdd m1_28490_22513# m1_28490_22513# m1_28090_22402# m1_28624_21786# m1_28624_21786#
+ pfet$183
Xpfet$183_21 vdd vdd vdd m1_21056_22402# m1_19839_21786# m1_19839_21786# pfet$183
Xpfet$190_2 vdd vdd m1_n789_25858# m1_326_24346# pfet$190
Xpfet$205_5 vdd vdd m1_n10308_24542# m1_n9952_24224# pfet$205
Xpfet$183_1 vdd m1_7388_22513# m1_7388_22513# m1_6988_22402# m1_7522_21786# m1_7522_21786#
+ pfet$183
Xpfet$183_10 vdd m1_3871_22513# m1_3871_22513# m1_2843_22102# m1_4637_21786# m1_4637_21786#
+ pfet$183
Xnfet$204_0 pd1 vss m1_n1263_21786# vss nfet$204
Xpfet$203_2 vdd m1_n4362_24346# m1_n4847_25662# m1_n4464_25980# pfet$203
Xnfet$201_12 m1_28470_16080# vss m1_28113_15778# vss nfet$201
Xpfet$181_102 vdd m1_28371_23922# m1_28635_24542# m1_28010_25858# pfet$181
Xnfet$198_15 m1_28624_21786# vss m1_29256_21786# vss nfet$198
Xnfet$195_7 m1_5771_21786# m1_5771_21786# m1_7388_22513# m1_7388_22513# m1_6992_21586#
+ vss nfet$195
Xpfet$187_8 vdd vdd m1_n1133_19550# m1_n7383_17599# pfet$187
Xpfet$186_10 vdd vdd m1_27031_17343# m1_n10452_25858# pfet$186
Xnfet$193_4 m1_12259_24224# m1_12259_24224# m1_11903_24542# m1_11903_24542# m1_12357_24542#
+ vss nfet$193
Xpfet$207_9 vdd vdd m1_n4464_25980# m1_n4623_25487# pfet$207
Xpfet$192_6 vdd vdd m1_31535_19792# m1_14422_22513# pfet$192
Xpfet$185_5 vdd vdd m1_1120_21786# m1_488_21786# pfet$185
Xnfet$195_16 m1_27003_21590# m1_27003_21590# m1_28490_22513# m1_28490_22513# m1_27462_21586#
+ vss nfet$195
Xnfet$213_5 m1_9944_16080# m1_9944_16080# m1_9485_17714# m1_9485_17714# m1_10042_16398#
+ vss nfet$213
Xnfet$220_6 m1_n5764_21786# m1_n5764_21786# vss vss m1_n6282_21430# vss nfet$220
Xnfet$206_4 m1_1120_21786# m1_1120_21786# vss vss m1_n42_21586# vss nfet$206
Xpfet$190_3 vdd m1_n646_24542# vdd m1_326_24346# pfet$190
Xpfet$205_6 vdd m1_n10308_24542# vdd m1_n9336_24346# pfet$205
Xpfet$183_2 vdd m1_7388_22513# m1_7388_22513# m1_6360_22102# m1_8154_21786# m1_8154_21786#
+ pfet$183
Xpfet$183_33 vdd m1_28490_22513# m1_28490_22513# m1_27462_22102# m1_29256_21786# m1_29256_21786#
+ pfet$183
Xpfet$183_22 vdd m1_21456_22513# m1_21456_22513# m1_20428_22102# m1_22222_21786# m1_22222_21786#
+ pfet$183
Xpfet$183_11 vdd vdd vdd m1_2843_22102# m1_2384_21590# m1_2384_21590# pfet$183
Xnfet$204_1 pd2 vss m1_2254_21786# vss nfet$204
Xpfet$203_3 vdd m1_n3184_24224# m1_n3651_26174# m1_n4623_25487# pfet$203
Xnfet$201_13 m1_26217_17714# vss m1_25747_17714# vss nfet$201
Xpfet$189_10 vdd vdd m1_35071_24542# m1_32675_25947# pfet$189
Xpfet$201_0 vdd vdd m1_n7513_20152# m1_35837_22102# pfet$201
Xpfet$181_103 vdd vdd m1_28635_24542# m1_28991_24224# pfet$181
Xnfet$195_8 m1_23486_21590# m1_23486_21590# m1_24973_22513# m1_24973_22513# m1_23945_21586#
+ vss nfet$195
Xnfet$198_16 m1_26873_21786# vss m1_27003_21590# vss nfet$198
Xpfet$187_9 vdd vdd m1_27003_19550# m1_25747_17714# pfet$187
Xpfet$186_11 vdd vdd m1_26807_17518# m1_26217_17714# pfet$186
Xpfet$199_0 vdd vdd m1_n7247_17714# m1_n6788_16080# pfet$199
Xnfet$193_5 m1_8692_24346# m1_8692_24346# vss vss m1_8174_24542# vss nfet$193
Xpfet$192_7 vdd vdd m1_31535_22102# m1_354_22513# pfet$192
Xnfet$227_0 m1_n927_19404# m1_n927_19404# vss vss m1_n6282_20470# vss nfet$227
Xpfet$185_6 vdd vdd m1_5901_21590# m1_5771_21786# pfet$185
Xnfet$195_17 m1_12935_21590# m1_12935_21590# m1_14422_22513# m1_14422_22513# m1_13394_21586#
+ vss nfet$195
Xnfet$213_6 m1_1578_16080# m1_1578_16080# vss vss m1_3141_17358# vss nfet$213
Xnfet$220_7 m1_n3822_21786# m1_n3822_21786# m1_n4485_21904# m1_n4485_21904# m1_n3724_21430#
+ vss nfet$220
Xnfet$206_5 m1_4005_21786# m1_4005_21786# vss vss m1_2843_21586# vss nfet$206
Xpfet$190_4 vdd vdd m1_32675_25947# m1_33790_24346# pfet$190
Xpfet$205_7 vdd vdd m1_n10452_25858# m1_n4978_24224# pfet$205
Xpfet$183_3 vdd m1_9645_21447# m1_9645_21447# m1_10505_22402# m1_11039_21786# m1_11039_21786#
+ pfet$183
Xpfet$183_34 vdd vdd vdd m1_28090_22402# m1_26873_21786# m1_26873_21786# pfet$183
Xpfet$183_23 vdd vdd vdd m1_23945_22102# m1_23486_21590# m1_23486_21590# pfet$183
Xpfet$183_12 vdd vdd vdd m1_3471_22402# m1_2254_21786# m1_2254_21786# pfet$183
Xnfet$204_2 pd9 vss m1_26873_21786# vss nfet$204
Xpfet$203_4 vdd m1_n2567_23922# m1_n3184_24224# m1_n4464_25980# pfet$203
Xpfet$181_0 vdd vdd m1_3049_25662# m1_2912_25858# pfet$181
Xpfet$189_11 vdd vdd m1_32817_25662# m1_32675_25947# pfet$189
Xpfet$181_104 vdd m1_25912_25658# m1_26705_24542# m1_23964_25662# pfet$181
Xnfet$198_17 m1_25107_21786# vss m1_25739_21786# vss nfet$198
Xnfet$195_9 m1_23356_21786# m1_23356_21786# m1_24973_22513# m1_24973_22513# m1_24577_21586#
+ vss nfet$195
Xpfet$186_12 vdd vdd m1_26676_16080# m1_n7513_20152# pfet$186
Xpfet$199_1 vdd m1_n7247_17714# vdd m1_n6172_16202# pfet$199
Xnfet$193_6 m1_8076_24224# m1_8076_24224# m1_7720_24542# m1_7720_24542# m1_8174_24542#
+ vss nfet$193
Xnfet$227_1 m1_n2543_20130# m1_n2543_20130# m1_n5227_20152# m1_n5227_20152# m1_n2445_20470#
+ vss nfet$227
Xpfet$185_7 vdd vdd m1_4637_21786# m1_4005_21786# pfet$185
Xnfet$213_7 m1_5761_16080# m1_5761_16080# m1_5302_17714# m1_5302_17714# m1_5859_16398#
+ vss nfet$213
Xnfet$220_8 m1_9624_19404# m1_9624_19404# vss vss m1_n3724_21430# vss nfet$220
Xnfet$206_6 m1_4637_21786# m1_4637_21786# vss vss m1_3475_21586# vss nfet$206
Xpfet$183_35 vdd vdd vdd m1_13394_22102# m1_12935_21590# m1_12935_21590# pfet$183
Xpfet$190_5 vdd m1_32675_25947# vdd m1_34278_25658# pfet$190
Xpfet$183_24 vdd m1_17939_22513# m1_17939_22513# m1_16911_22102# m1_18705_21786# m1_18705_21786#
+ pfet$183
Xpfet$183_13 vdd vdd vdd m1_6988_22402# m1_5771_21786# m1_5771_21786# pfet$183
Xpfet$183_4 vdd vdd vdd m1_9877_22102# m1_9418_21590# m1_9418_21590# pfet$183
Xpfet$181_1 vdd m1_3536_25662# m1_3273_23922# m1_3049_25662# pfet$181
Xpfet$203_5 vdd m1_n10572_23922# m1_n10308_24542# m1_n10933_25858# pfet$203
Xnfet$202_0 m1_n10452_25858# vss m1_n1271_25858# vss nfet$202
Xpfet$189_12 vdd vdd m1_32193_25858# m1_25107_21786# pfet$189
Xpfet$181_105 vdd vdd m1_30888_24542# m1_28492_25858# pfet$181
Xpfet$181_90 vdd vdd m1_24309_25858# m1_25424_24346# pfet$181
Xpfet$199_2 vdd vdd m1_n5461_18030# m1_n5351_15778# pfet$199
Xpfet$186_13 vdd vdd m1_25747_17714# m1_26217_17714# pfet$186
Xnfet$193_7 m1_9180_25658# m1_9180_25658# vss vss m1_9639_25502# vss nfet$193
Xpfet$185_8 vdd vdd m1_2384_21590# m1_2254_21786# pfet$185
Xnfet$206_7 m1_488_21786# m1_488_21786# vss vss m1_n674_21586# vss nfet$206
Xnfet$213_8 m1_3015_15778# m1_3015_15778# m1_2905_18030# m1_2905_18030# m1_3141_17358#
+ vss nfet$213
Xnfet$220_9 m1_n6380_21786# m1_n6380_21786# m1_n6839_21786# m1_n6839_21786# m1_n6282_21430#
+ vss nfet$220
Xpfet$190_6 vdd vdd m1_32818_24542# m1_33174_24224# pfet$190
Xpfet$183_25 vdd m1_17939_22513# m1_17939_22513# m1_17539_22402# m1_18073_21786# m1_18073_21786#
+ pfet$183
Xpfet$183_14 vdd vdd vdd m1_n46_22402# m1_n1263_21786# m1_n1263_21786# pfet$183
Xpfet$183_5 vdd m1_9645_21447# m1_9645_21447# m1_9877_22102# m1_11671_21786# m1_11671_21786#
+ pfet$183
Xpfet$181_2 vdd vdd m1_3394_25858# m1_4509_24346# pfet$181
Xpfet$203_6 vdd m1_n8848_25658# m1_n8055_24542# m1_n10796_25662# pfet$203
Xnfet$202_1 m1_n789_25858# vss m1_n647_25662# vss nfet$202
Xpfet$189_13 vdd vdd m1_33790_24346# m1_n7513_20152# pfet$189
Xpfet$181_106 vdd vdd m1_25107_21786# m1_28492_25858# pfet$181
Xpfet$181_91 vdd vdd m1_23356_21786# pd8 pfet$181
Xpfet$181_80 vdd vdd m1_17058_24346# m1_n7513_20152# pfet$181
Xpfet$199_3 vdd m1_n5461_18030# vdd m1_n6788_16080# pfet$199
Xpfet$185_9 vdd vdd m1_22222_21786# m1_21590_21786# pfet$185
Xnfet$193_8 m1_8692_24346# m1_8692_24346# m1_7577_25858# m1_7577_25858# m1_9639_25502#
+ vss nfet$193
Xpfet$197_0 vdd vdd fout m1_34093_22102# pfet$197
Xnfet$206_8 m1_25739_21786# m1_25739_21786# vss vss m1_24577_21586# vss nfet$206
Xnfet$213_9 m1_2194_16202# m1_2194_16202# vss vss m1_1676_16398# vss nfet$213
Xpfet$190_7 vdd m1_32818_24542# vdd m1_33790_24346# pfet$190
Xpfet$183_26 vdd vdd vdd m1_16911_22102# m1_16452_21590# m1_16452_21590# pfet$183
Xpfet$183_15 vdd m1_354_22513# m1_354_22513# m1_n46_22402# m1_488_21786# m1_488_21786#
+ pfet$183
Xnfet$225_0 m1_n8283_20611# vss m1_n8283_19850# vss nfet$225
Xpfet$183_6 vdd vdd vdd m1_10505_22402# m1_9288_21786# m1_9288_21786# pfet$183
Xpfet$203_7 vdd m1_n3541_23922# m1_n4362_24346# m1_n4623_25487# pfet$203
Xpfet$181_3 vdd m1_3394_25858# vdd m1_4997_25658# pfet$181
Xnfet$202_2 m1_n1271_25858# vss m1_n1134_25662# vss nfet$202
Xpfet$181_107 vdd m1_24309_25858# vdd m1_25912_25658# pfet$181
Xnfet$193_20 m1_21241_24346# m1_21241_24346# m1_20126_25858# m1_20126_25858# m1_22188_25502#
+ vss nfet$193
Xpfet$181_92 vdd vdd m1_28492_25858# m1_29607_24346# pfet$181
Xpfet$181_81 vdd vdd m1_18339_24542# m1_15943_25858# pfet$181
Xpfet$181_70 vdd vdd m1_14156_24542# m1_11760_25858# pfet$181
Xpfet$199_4 vdd vdd m1_26217_17714# m1_26676_16080# pfet$199
Xnfet$193_9 m1_17058_24346# m1_17058_24346# vss vss m1_16540_24542# vss nfet$193
Xnfet$206_9 m1_25107_21786# m1_25107_21786# vss vss m1_23945_21586# vss nfet$206
Xnfet$225_1 m1_n7513_20152# m1_n8283_19850# vss vss nfet$225
Xnfet$218_0 m1_n10452_25858# m1_n10452_25858# m1_n7186_25858# m1_n7186_25858# m1_n6629_25502#
+ vss nfet$218
Xpfet$183_7 vdd m1_354_22513# m1_354_22513# m1_n674_22102# m1_1120_21786# m1_1120_21786#
+ pfet$183
Xpfet$183_27 vdd m1_14422_22513# m1_14422_22513# m1_14022_22402# m1_14556_21786# m1_14556_21786#
+ pfet$183
Xpfet$183_16 vdd m1_24973_22513# m1_24973_22513# m1_23945_22102# m1_25739_21786# m1_25739_21786#
+ pfet$183
Xpfet$181_4 vdd vdd m1_3893_24224# m1_3273_23922# pfet$181
Xnfet$202_3 m1_n7513_20152# vss m1_326_24346# vss nfet$202
Xpfet$181_108 vdd vdd m1_25424_24346# m1_n7513_20152# pfet$181
Xnfet$193_21 m1_28991_24224# m1_28991_24224# m1_28635_24542# m1_28635_24542# m1_29089_24542#
+ vss nfet$193
Xnfet$193_10 m1_17546_25658# m1_17546_25658# vss vss m1_18005_25502# vss nfet$193
Xnfet$200_0 sd9 vss m1_n7401_15478# vss nfet$200
Xpfet$181_93 vdd m1_28991_24224# m1_30095_25658# m1_28010_25858# pfet$181
Xpfet$181_82 vdd vdd m1_21241_24346# m1_n7513_20152# pfet$181
Xpfet$181_71 vdd vdd m1_11039_21786# m1_11760_25858# pfet$181
Xpfet$181_60 vdd vdd m1_20126_25858# m1_21241_24346# pfet$181
Xpfet$199_5 vdd m1_26217_17714# vdd m1_27292_16202# pfet$199
Xnfet$198_0 m1_n1263_21786# vss m1_n1133_21590# vss nfet$198
Xnfet$225_2 m1_n8145_21908# vss m1_n8283_20611# vss nfet$225
Xnfet$218_1 m1_n6111_25858# m1_n6111_25858# vss vss m1_n6629_25502# vss nfet$218
Xpfet$183_8 vdd vdd vdd m1_6360_22102# m1_5901_21590# m1_5901_21590# pfet$183
Xpfet$183_28 vdd m1_14422_22513# m1_14422_22513# m1_13394_22102# m1_15188_21786# m1_15188_21786#
+ pfet$183
Xpfet$183_17 vdd m1_21456_22513# m1_21456_22513# m1_21056_22402# m1_21590_21786# m1_21590_21786#
+ pfet$183
Xnfet$196_10 m1_9015_17714# m1_9015_17714# vss vss m1_14005_20470# vss nfet$196
Xpfet$181_5 vdd m1_3893_24224# m1_4997_25658# m1_2912_25858# pfet$181
Xnfet$202_4 m1_n789_25858# vss m1_1607_24542# vss nfet$202
Xpfet$181_109 vdd m1_12259_24224# m1_13363_25658# m1_11278_25858# pfet$181
Xnfet$193_22 m1_29607_24346# m1_29607_24346# vss vss m1_29089_24542# vss nfet$193
Xnfet$193_11 m1_16442_24224# m1_16442_24224# m1_16086_24542# m1_16086_24542# m1_16540_24542#
+ vss nfet$193
Xnfet$200_1 sd2 vss m1_21880_15478# vss nfet$200
Xpfet$181_94 vdd m1_28492_25858# vdd m1_30095_25658# pfet$181
Xpfet$181_83 vdd m1_21729_25658# m1_22522_24542# m1_19781_25662# pfet$181
Xpfet$181_72 vdd m1_13363_25658# m1_14156_24542# m1_11415_25662# pfet$181
Xpfet$181_61 vdd m1_24452_24542# vdd m1_25424_24346# pfet$181
Xpfet$181_50 vdd vdd m1_20268_25662# m1_20126_25858# pfet$181
Xpfet$199_6 vdd vdd m1_28003_18030# m1_28113_15778# pfet$199
Xnfet$199_10 m1_26063_15478# vss m1_29239_20152# vss nfet$199
Xnfet$198_1 m1_11039_21786# vss m1_11671_21786# vss nfet$198
Xnfet$225_3 m1_n8283_19850# m1_n8283_20611# vss vss nfet$225
Xpfet$195_0 vdd m1_34093_22102# vdd m1_28490_22513# pfet$195
Xpfet$183_29 vdd vdd vdd m1_14022_22402# m1_12805_21786# m1_12805_21786# pfet$183
Xpfet$183_18 vdd vdd vdd m1_24573_22402# m1_23356_21786# m1_23356_21786# pfet$183
Xpfet$183_9 vdd m1_3871_22513# m1_3871_22513# m1_3471_22402# m1_4005_21786# m1_4005_21786#
+ pfet$183
Xnfet$196_11 m1_13198_17714# m1_13198_17714# vss vss m1_17522_20470# vss nfet$196
Xpfet$181_6 vdd vdd m1_3536_25662# m1_3394_25858# pfet$181
Xnfet$223_0 m1_n10933_25858# m1_n8848_25658# m1_n8055_24542# vss nfet$223
Xpfet$208_0 vdd vdd m1_n7186_25858# m1_n10452_25858# pfet$208
Xnfet$202_5 m1_n789_25858# vss m1_488_21786# vss nfet$202
Xnfet$200_2 sd1 vss m1_26063_15478# vss nfet$200
Xnfet$193_23 m1_25424_24346# m1_25424_24346# m1_24309_25858# m1_24309_25858# m1_26371_25502#
+ vss nfet$193
Xnfet$193_12 m1_17058_24346# m1_17058_24346# m1_15943_25858# m1_15943_25858# m1_18005_25502#
+ vss nfet$193
Xpfet$181_95 vdd vdd m1_28991_24224# m1_28371_23922# pfet$181
Xpfet$181_84 vdd vdd m1_23827_25858# m1_18073_21786# pfet$181
Xpfet$181_73 vdd m1_16086_24542# vdd m1_17058_24346# pfet$181
Xpfet$181_62 vdd vdd m1_24452_24542# m1_24808_24224# pfet$181
Xpfet$181_51 vdd vdd m1_20625_24224# m1_20005_23922# pfet$181
Xpfet$181_40 vdd vdd m1_11760_25858# m1_12875_24346# pfet$181
Xpfet$199_7 vdd m1_28003_18030# vdd m1_26676_16080# pfet$199
Xnfet$199_11 m1_9331_15478# vss m1_15171_20152# vss nfet$199
Xnfet$198_2 m1_12805_21786# vss m1_12935_21590# vss nfet$198
Xpfet$183_19 vdd m1_24973_22513# m1_24973_22513# m1_24573_22402# m1_25107_21786# m1_25107_21786#
+ pfet$183
Xpfet$195_1 vdd vdd m1_34093_22102# m1_34843_21786# pfet$195
Xpfet$188_0 vdd vdd m1_n7401_15478# sd9 pfet$188
Xnfet$196_12 m1_16452_19550# m1_16452_19550# vss vss m1_16890_20470# vss nfet$196
Xpfet$181_7 vdd vdd m1_7232_25662# m1_7095_25858# pfet$181
Xnfet$216_0 m1_n6274_17836# m1_n4994_16080# m1_n5461_18030# vss nfet$216
Xnfet$223_1 m1_n10796_25662# m1_n10572_23922# m1_n10308_24542# vss nfet$223
Xpfet$208_1 vdd m1_n7186_25858# vdd m1_n6111_25858# pfet$208
Xnfet$202_6 m1_n910_23922# vss m1_n290_24224# vss nfet$202
Xnfet$193_24 m1_30095_25658# m1_30095_25658# vss vss m1_30554_25502# vss nfet$193
Xnfet$193_13 m1_13363_25658# m1_13363_25658# vss vss m1_13822_25502# vss nfet$193
Xpfet$181_96 vdd m1_28635_24542# vdd m1_29607_24346# pfet$181
Xpfet$181_85 vdd m1_24188_23922# m1_24452_24542# m1_23827_25858# pfet$181
Xpfet$181_74 vdd vdd m1_14556_21786# m1_15943_25858# pfet$181
Xpfet$181_63 vdd vdd m1_19781_25662# m1_19644_25858# pfet$181
Xpfet$181_52 vdd m1_20268_25662# m1_20005_23922# m1_19781_25662# pfet$181
Xpfet$181_41 vdd vdd m1_9288_21786# pd4 pfet$181
Xpfet$181_30 vdd vdd m1_2912_25858# m1_488_21786# pfet$181
Xnfet$199_12 m1_13514_15478# vss m1_18688_20152# vss nfet$199
Xnfet$198_3 m1_9288_21786# vss m1_9418_21590# vss nfet$198
Xnfet$196_0 m1_n3534_17714# m1_n3534_17714# vss vss m1_3454_20470# vss nfet$196
Xpfet$195_2 vdd vdd m1_30256_22102# m1_7388_22513# pfet$195
Xpfet$188_1 vdd vdd m1_21880_15478# sd2 pfet$188
Xnfet$196_13 m1_19969_19550# m1_19969_19550# vss vss m1_20407_20470# vss nfet$196
Xnfet$223_2 m1_n10933_25858# m1_n10309_25662# m1_n10572_23922# vss nfet$223
Xnfet$209_0 m1_31535_22102# m1_32818_21586# vss vss nfet$209
Xpfet$181_8 vdd vdd m1_8076_24224# m1_7456_23922# pfet$181
Xnfet$216_1 m1_n6433_17343# m1_n4377_15778# m1_n4994_16080# vss nfet$216
Xnfet$202_7 m1_25107_21786# vss m1_32193_25858# vss nfet$202
Xpfet$184_30 vdd vdd vdd m1_24560_19550# m1_21880_15478# m1_21880_15478# pfet$184
Xpfet$213_0 vdd vdd m1_n8145_21908# m1_n6839_20152# pfet$213
Xnfet$193_25 m1_29607_24346# m1_29607_24346# m1_28492_25858# m1_28492_25858# m1_30554_25502#
+ vss nfet$193
Xnfet$193_14 m1_12875_24346# m1_12875_24346# m1_11760_25858# m1_11760_25858# m1_13822_25502#
+ vss nfet$193
Xnfet$202_10 m1_32675_25947# vss m1_35071_24542# vss nfet$202
Xpfet$181_97 vdd vdd m1_21590_21786# m1_24309_25858# pfet$181
Xpfet$181_86 vdd m1_28634_25662# m1_28371_23922# m1_28147_25662# pfet$181
Xpfet$181_75 vdd vdd m1_19644_25858# m1_14556_21786# pfet$181
Xpfet$181_64 vdd vdd m1_22522_24542# m1_20126_25858# pfet$181
Xpfet$181_53 vdd m1_20625_24224# m1_21729_25658# m1_19644_25858# pfet$181
Xpfet$181_42 vdd m1_11760_25858# vdd m1_13363_25658# pfet$181
Xpfet$181_31 vdd m1_3273_23922# m1_3537_24542# m1_2912_25858# pfet$181
Xpfet$181_20 vdd vdd m1_4509_24346# m1_n7513_20152# pfet$181
Xnfet$213_20 m1_22493_16080# m1_22493_16080# m1_22034_17714# m1_22034_17714# m1_22591_16398#
+ vss nfet$213
Xnfet$199_13 m1_13198_17714# vss m1_16452_19550# vss nfet$199
Xnfet$198_4 m1_7522_21786# vss m1_8154_21786# vss nfet$198
Xnfet$196_1 m1_2384_19550# m1_2384_19550# vss vss m1_2822_20470# vss nfet$196
Xpfet$188_2 vdd vdd m1_26063_15478# sd1 pfet$188
Xpfet$195_3 vdd m1_31535_22102# vdd m1_3871_22513# pfet$195
Xnfet$196_14 m1_17381_17714# m1_17381_17714# vss vss m1_21039_20470# vss nfet$196
Xpfet$181_9 vdd m1_7719_25662# m1_7456_23922# m1_7232_25662# pfet$181
Xnfet$216_2 m1_n6274_17836# m1_n5351_15778# m1_n6172_16202# vss nfet$216
Xnfet$223_3 m1_n10796_25662# m1_n9952_24224# m1_n8848_25658# vss nfet$223
Xpfet$184_31 vdd m1_n2543_20130# m1_n2543_20130# m1_20407_19850# m1_19969_19550# m1_19969_19550#
+ pfet$184
Xpfet$184_20 vdd m1_n3822_21786# m1_n3822_21786# m1_14009_19550# m1_9015_17714# m1_9015_17714#
+ pfet$184
Xpfet$193_0 vdd m1_n647_25662# m1_n910_23922# m1_n1134_25662# pfet$193
Xnfet$202_8 m1_32193_25858# vss m1_32330_25662# vss nfet$202
Xnfet$221_0 m1_n8625_26174# vss m1_n8055_24542# vss nfet$221
Xpfet$206_0 vdd vdd m1_n4485_20152# m1_n3822_20130# pfet$206
Xnfet$193_26 m1_25912_25658# m1_25912_25658# vss vss m1_26371_25502# vss nfet$193
Xnfet$193_15 m1_25424_24346# m1_25424_24346# vss vss m1_24906_24542# vss nfet$193
Xnfet$202_11 m1_32554_23922# vss m1_33174_24224# vss nfet$202
Xpfet$181_98 vdd m1_30095_25658# m1_30888_24542# m1_28147_25662# pfet$181
Xpfet$181_87 vdd vdd m1_28147_25662# m1_28010_25858# pfet$181
Xpfet$181_76 vdd m1_20005_23922# m1_20269_24542# m1_19644_25858# pfet$181
Xpfet$181_65 vdd vdd m1_18073_21786# m1_20126_25858# pfet$181
Xpfet$181_54 vdd vdd m1_24808_24224# m1_24188_23922# pfet$181
Xpfet$181_43 vdd vdd m1_12805_21786# pd5 pfet$181
Xpfet$181_32 vdd vdd m1_7720_24542# m1_8076_24224# pfet$181
Xpfet$181_21 vdd m1_7456_23922# m1_7720_24542# m1_7095_25858# pfet$181
Xpfet$181_10 vdd m1_8076_24224# m1_9180_25658# m1_7095_25858# pfet$181
Xnfet$194_80 m1_28147_25662# m1_28991_24224# m1_30095_25658# vss nfet$194
Xnfet$213_21 m1_14127_16080# m1_14127_16080# vss vss m1_15690_17358# vss nfet$213
Xnfet$213_10 m1_1578_16080# m1_1578_16080# m1_1119_17714# m1_1119_17714# m1_1676_16398#
+ vss nfet$213
Xnfet$199_14 m1_21564_17714# vss m1_23486_19550# vss nfet$199
Xnfet$198_5 m1_488_21786# vss m1_1120_21786# vss nfet$198
Xpfet$195_4 vdd m1_30256_22102# vdd m1_9645_21447# pfet$195
Xnfet$196_2 m1_5901_19550# m1_5901_19550# vss vss m1_6339_20470# vss nfet$196
Xnfet$196_15 m1_21564_17714# m1_21564_17714# vss vss m1_24556_20470# vss nfet$196
Xnfet$216_3 m1_n6433_17343# m1_n6172_16202# m1_n6657_17518# vss nfet$216
Xnfet$223_4 m1_n4623_25487# m1_n2567_23922# m1_n3184_24224# vss nfet$223
Xpfet$184_32 vdd m1_n2543_20130# m1_n2543_20130# m1_21043_19550# m1_17381_17714# m1_17381_17714#
+ pfet$184
Xpfet$184_21 vdd vdd vdd m1_13373_19850# m1_15171_20152# m1_15171_20152# pfet$184
Xpfet$184_10 vdd vdd vdd m1_9856_19850# m1_11654_20152# m1_11654_20152# pfet$184
Xpfet$186_0 vdd vdd m1_n6274_17836# m1_n6433_17343# pfet$186
Xnfet$221_10 vss vss m1_n4978_24224# vss nfet$221
Xpfet$193_1 vdd m1_n910_23922# m1_n646_24542# m1_n1271_25858# pfet$193
Xnfet$202_9 m1_n7513_20152# vss m1_33790_24346# vss nfet$202
Xnfet$197_80 m1_18824_17836# m1_19747_15778# m1_18926_16202# vss nfet$197
Xnfet$214_0 m1_4620_20152# m1_4620_20152# m1_2590_19404# m1_2590_19404# m1_3454_20470#
+ vss nfet$214
Xpfet$206_1 vdd m1_n4485_21904# vdd m1_9624_19404# pfet$206
Xnfet$221_1 m1_n8625_26174# vss m1_n7082_23622# vss nfet$221
Xnfet$193_27 m1_12875_24346# m1_12875_24346# vss vss m1_12357_24542# vss nfet$193
Xnfet$193_16 m1_24808_24224# m1_24808_24224# m1_24452_24542# m1_24452_24542# m1_24906_24542#
+ vss nfet$193
Xpfet$181_99 vdd vdd m1_26705_24542# m1_24309_25858# pfet$181
Xnfet$202_12 m1_32675_25947# vss m1_28624_21786# vss nfet$202
Xpfet$181_88 vdd vdd m1_28634_25662# m1_28492_25858# pfet$181
Xpfet$181_77 vdd vdd m1_20269_24542# m1_20625_24224# pfet$181
Xpfet$181_66 vdd vdd m1_15461_25858# m1_11039_21786# pfet$181
Xpfet$181_55 vdd m1_24451_25662# m1_24188_23922# m1_23964_25662# pfet$181
Xpfet$181_44 vdd m1_15943_25858# vdd m1_17546_25658# pfet$181
Xpfet$181_33 vdd vdd m1_7522_21786# m1_7577_25858# pfet$181
Xpfet$181_22 vdd vdd m1_3537_24542# m1_3893_24224# pfet$181
Xpfet$181_11 vdd vdd m1_7719_25662# m1_7577_25858# pfet$181
Xnfet$194_81 m1_n7513_20152# vss m1_25424_24346# vss nfet$194
Xnfet$194_70 m1_21590_21786# vss m1_28010_25858# vss nfet$194
Xnfet$213_22 m1_15564_15778# m1_15564_15778# m1_15454_18030# m1_15454_18030# m1_15690_17358#
+ vss nfet$213
Xnfet$213_11 m1_6377_16202# m1_6377_16202# vss vss m1_5859_16398# vss nfet$213
Xnfet$199_15 m1_17697_15478# vss m1_22205_20152# vss nfet$199
Xnfet$198_6 m1_5771_21786# vss m1_5901_21590# vss nfet$198
Xpfet$187_10 vdd vdd m1_29239_20152# m1_26063_15478# pfet$187
Xnfet$196_3 m1_4832_17714# m1_4832_17714# vss vss m1_10488_20470# vss nfet$196
Xnfet$196_16 m1_23486_19550# m1_23486_19550# vss vss m1_23924_20470# vss nfet$196
Xnfet$216_4 m1_27031_17343# m1_27292_16202# m1_26807_17518# vss nfet$216
Xnfet$223_5 m1_n4464_25980# m1_n3541_23922# m1_n4362_24346# vss nfet$223
Xnfet$194_0 m1_3394_25858# vss m1_5790_24542# vss nfet$194
Xpfet$184_33 vdd m1_n3206_20274# m1_n3206_20274# m1_24560_19550# m1_21564_17714# m1_21564_17714#
+ pfet$184
Xpfet$184_22 vdd vdd vdd m1_14009_19550# m1_9331_15478# m1_9331_15478# pfet$184
Xpfet$184_11 vdd vdd vdd m1_10492_19550# m1_5148_15478# m1_5148_15478# pfet$184
Xpfet$186_1 vdd vdd m1_n4377_15778# m1_n7247_17714# pfet$186
Xnfet$221_11 m1_n10452_25858# vss m1_n4847_25662# vss nfet$221
Xpfet$193_2 vdd m1_n290_24224# m1_814_25658# m1_n1271_25858# pfet$193
Xnfet$197_81 m1_13198_17714# vss m1_10299_17343# vss nfet$197
Xnfet$197_70 m1_n7513_20152# vss m1_18310_16080# vss nfet$197
Xnfet$207_0 m1_21456_22513# m1_21456_22513# m1_30256_19792# m1_30256_19792# m1_30492_20470#
+ vss nfet$207
Xnfet$214_1 m1_1103_20152# m1_1103_20152# m1_n927_19404# m1_n927_19404# m1_n63_20470#
+ vss nfet$214
Xpfet$206_2 vdd m1_n5227_21418# vdd m1_2590_19404# pfet$206
Xnfet$221_2 vss vss m1_n9336_24346# vss nfet$221
Xnfet$193_17 m1_20625_24224# m1_20625_24224# m1_20269_24542# m1_20269_24542# m1_20723_24542#
+ vss nfet$193
Xnfet$202_13 m1_32675_25947# vss m1_32817_25662# vss nfet$202
Xpfet$181_89 vdd vdd m1_19839_21786# pd7 pfet$181
Xpfet$181_78 vdd m1_20269_24542# vdd m1_21241_24346# pfet$181
Xpfet$181_67 vdd m1_15822_23922# m1_16086_24542# m1_15461_25858# pfet$181
Xpfet$181_56 vdd m1_24808_24224# m1_25912_25658# m1_23827_25858# pfet$181
Xpfet$181_45 vdd vdd m1_16442_24224# m1_15822_23922# pfet$181
Xpfet$181_34 vdd m1_9180_25658# m1_9973_24542# m1_7232_25662# pfet$181
Xpfet$181_23 vdd m1_3537_24542# vdd m1_4509_24346# pfet$181
Xpfet$181_12 vdd m1_7577_25858# vdd m1_9180_25658# pfet$181
Xpfet$211_0 vdd vdd m1_n5227_20152# m1_n2543_20130# pfet$211
Xnfet$194_82 m1_11415_25662# m1_12259_24224# m1_13363_25658# vss nfet$194
Xnfet$194_71 m1_28147_25662# m1_28371_23922# m1_28635_24542# vss nfet$194
Xnfet$194_60 pd6 vss m1_16322_21786# vss nfet$194
Xnfet$213_23 m1_18926_16202# m1_18926_16202# vss vss m1_18408_16398# vss nfet$213
Xnfet$213_12 m1_n1168_15778# m1_n1168_15778# m1_n1278_18030# m1_n1278_18030# m1_n1042_17358#
+ vss nfet$213
Xnfet$199_16 m1_17381_17714# vss m1_19969_19550# vss nfet$199
Xnfet$198_7 m1_4005_21786# vss m1_4637_21786# vss nfet$198
Xpfet$187_11 vdd vdd m1_18688_20152# m1_13514_15478# pfet$187
Xnfet$196_4 m1_9418_19550# m1_9418_19550# vss vss m1_9856_20470# vss nfet$196
Xnfet$196_17 m1_12935_19550# m1_12935_19550# vss vss m1_13373_20470# vss nfet$196
Xnfet$216_5 m1_27031_17343# m1_29087_15778# m1_28470_16080# vss nfet$216
Xnfet$223_6 m1_n4464_25980# m1_n3184_24224# m1_n3651_26174# vss nfet$223
Xpfet$193_3 vdd m1_814_25658# m1_1607_24542# m1_n1134_25662# pfet$193
Xpfet$186_2 vdd vdd m1_n5351_15778# m1_n4994_16080# pfet$186
Xnfet$194_1 m1_2912_25858# m1_4997_25658# m1_5790_24542# vss nfet$194
Xpfet$184_34 vdd m1_n3206_20274# m1_n3206_20274# m1_23924_19850# m1_23486_19550# m1_23486_19550#
+ pfet$184
Xpfet$184_23 vdd vdd vdd m1_16890_19850# m1_18688_20152# m1_18688_20152# pfet$184
Xpfet$184_12 vdd m1_6107_19404# m1_6107_19404# m1_6975_19550# m1_649_17714# m1_649_17714#
+ pfet$184
Xnfet$221_12 m1_n10452_25858# vss m1_n5571_25662# vss nfet$221
Xnfet$207_1 m1_14422_22513# m1_14422_22513# m1_31535_19792# m1_31535_19792# m1_31771_20470#
+ vss nfet$207
Xnfet$214_2 m1_n3218_15478# m1_n3218_15478# m1_2590_19404# m1_2590_19404# m1_2822_20470#
+ vss nfet$214
Xnfet$221_3 fin vss m1_n10933_25858# vss nfet$221
Xnfet$197_82 m1_10299_17343# vss m1_10458_17836# vss nfet$197
Xpfet$191_0 vdd vdd vdd m1_33050_22344# m1_31535_22102# m1_31535_22102# pfet$191
Xnfet$197_71 m1_14641_17836# m1_15921_16080# m1_15454_18030# vss nfet$197
Xnfet$197_60 m1_18665_17343# vss m1_18824_17836# vss nfet$197
Xpfet$206_3 vdd vdd m1_n5227_21418# m1_6107_19404# pfet$206
Xnfet$193_18 m1_21241_24346# m1_21241_24346# vss vss m1_20723_24542# vss nfet$193
Xpfet$181_79 vdd m1_17546_25658# m1_18339_24542# m1_15598_25662# pfet$181
Xpfet$181_68 vdd vdd m1_16086_24542# m1_16442_24224# pfet$181
Xpfet$181_57 vdd vdd m1_24451_25662# m1_24309_25858# pfet$181
Xpfet$181_46 vdd m1_16442_24224# m1_17546_25658# m1_15461_25858# pfet$181
Xpfet$181_35 vdd m1_7720_24542# vdd m1_8692_24346# pfet$181
Xpfet$181_24 vdd vdd m1_5790_24542# m1_3394_25858# pfet$181
Xpfet$181_13 vdd vdd m1_12259_24224# m1_11639_23922# pfet$181
Xpfet$211_1 vdd m1_n4485_20152# vdd m1_n3206_20274# pfet$211
Xpfet$204_0 vdd vdd m1_n7320_25516# m1_n7186_25858# pfet$204
Xnfet$194_72 m1_23827_25858# m1_25912_25658# m1_26705_24542# vss nfet$194
Xnfet$194_61 m1_23964_25662# m1_24808_24224# m1_25912_25658# vss nfet$194
Xnfet$194_50 m1_n7513_20152# vss m1_21241_24346# vss nfet$194
Xnfet$213_24 m1_18310_16080# m1_18310_16080# m1_17851_17714# m1_17851_17714# m1_18408_16398#
+ vss nfet$213
Xnfet$213_13 m1_n2605_16080# m1_n2605_16080# vss vss m1_n1042_17358# vss nfet$213
Xnfet$199_17 m1_21880_15478# vss m1_25722_20152# vss nfet$199
Xnfet$198_8 m1_2254_21786# vss m1_2384_21590# vss nfet$198
Xpfet$187_12 vdd vdd m1_15171_20152# m1_9331_15478# pfet$187
Xnfet$196_5 m1_649_17714# m1_649_17714# vss vss m1_6971_20470# vss nfet$196
Xnfet$223_7 m1_n4623_25487# m1_n4362_24346# m1_n4847_25662# vss nfet$223
Xpfet$193_4 vdd m1_33174_24224# m1_34278_25658# m1_32193_25858# pfet$193
Xnfet$216_6 m1_27190_17836# m1_28113_15778# m1_27292_16202# vss nfet$216
Xnfet$194_2 m1_n7513_20152# vss m1_4509_24346# vss nfet$194
Xpfet$184_35 vdd m1_n3822_21786# m1_n3822_21786# m1_13373_19850# m1_12935_19550# m1_12935_19550#
+ pfet$184
Xpfet$184_24 vdd m1_n1927_20274# m1_n1927_20274# m1_16890_19850# m1_16452_19550# m1_16452_19550#
+ pfet$184
Xpfet$184_13 vdd m1_n927_19404# m1_n927_19404# m1_n695_19850# m1_n1133_19550# m1_n1133_19550#
+ pfet$184
Xpfet$186_3 vdd vdd m1_n6657_17518# m1_n7247_17714# pfet$186
Xnfet$221_13 fin vss m1_n4623_25487# vss nfet$221
Xnfet$207_2 m1_17939_22513# m1_17939_22513# vss vss m1_31771_20470# vss nfet$207
Xnfet$214_3 m1_8137_20152# m1_8137_20152# m1_6107_19404# m1_6107_19404# m1_6971_20470#
+ vss nfet$214
Xnfet$221_4 m1_n10572_23922# vss m1_n9952_24224# vss nfet$221
Xnfet$197_72 m1_17851_17714# vss m1_18441_17518# vss nfet$197
Xnfet$197_61 m1_20104_16080# vss m1_19747_15778# vss nfet$197
Xnfet$197_50 m1_25747_17714# vss m1_22848_17343# vss nfet$197
Xpfet$184_0 vdd m1_2590_19404# m1_2590_19404# m1_3458_19550# m1_n3534_17714# m1_n3534_17714#
+ pfet$184
Xpfet$206_4 vdd vdd m1_n4485_21904# m1_n3822_21786# pfet$206
Xnfet$193_19 m1_21729_25658# m1_21729_25658# vss vss m1_22188_25502# vss nfet$193
Xnfet$212_0 fout vss m1_35837_22102# vss nfet$212
Xpfet$181_14 vdd vdd m1_11902_25662# m1_11760_25858# pfet$181
Xpfet$211_2 vdd m1_n5227_20152# vdd m1_n1927_20274# pfet$211
Xpfet$181_69 vdd vdd m1_12875_24346# m1_n7513_20152# pfet$181
Xpfet$181_58 vdd vdd m1_23964_25662# m1_23827_25858# pfet$181
Xpfet$181_47 vdd vdd m1_15943_25858# m1_17058_24346# pfet$181
Xpfet$181_36 vdd vdd m1_8692_24346# m1_n7513_20152# pfet$181
Xpfet$181_25 vdd vdd m1_4005_21786# m1_3394_25858# pfet$181
Xpfet$204_1 vdd vdd m1_n6111_25858# m1_n6856_24542# pfet$204
Xnfet$194_73 m1_24309_25858# vss m1_21590_21786# vss nfet$194
Xnfet$194_62 m1_24188_23922# vss m1_24808_24224# vss nfet$194
Xnfet$194_51 m1_19644_25858# m1_21729_25658# m1_22522_24542# vss nfet$194
Xnfet$194_40 m1_15598_25662# m1_16442_24224# m1_17546_25658# vss nfet$194
Xnfet$213_25 m1_14743_16202# m1_14743_16202# vss vss m1_14225_16398# vss nfet$213
Xnfet$213_14 m1_n2605_16080# m1_n2605_16080# m1_n3064_17714# m1_n3064_17714# m1_n2507_16398#
+ vss nfet$213
Xnfet$198_9 m1_23356_21786# vss m1_23486_21590# vss nfet$198
Xpfet$182_90 vdd m1_19747_15778# m1_18926_16202# m1_18665_17343# pfet$182
Xpfet$187_13 vdd vdd m1_16452_19550# m1_13198_17714# pfet$187
Xnfet$196_6 m1_n1133_19550# m1_n1133_19550# vss vss m1_n695_20470# vss nfet$196
Xnfet$216_7 m1_27190_17836# m1_28470_16080# m1_28003_18030# vss nfet$216
Xnfet$194_3 m1_488_21786# vss m1_2912_25858# vss nfet$194
Xpfet$193_5 vdd m1_32817_25662# m1_32554_23922# m1_32330_25662# pfet$193
Xpfet$184_25 vdd vdd vdd m1_17526_19550# m1_13514_15478# m1_13514_15478# pfet$184
Xpfet$184_14 vdd m1_n927_19404# m1_n927_19404# m1_n59_19550# m1_n7383_17599# m1_n7383_17599#
+ pfet$184
Xpfet$186_4 vdd vdd m1_n6433_17343# m1_n3534_17714# pfet$186
Xnfet$207_3 m1_24973_22513# m1_24973_22513# vss vss m1_30492_20470# vss nfet$207
Xnfet$214_4 m1_965_15478# m1_965_15478# m1_6107_19404# m1_6107_19404# m1_6339_20470#
+ vss nfet$214
Xnfet$221_5 m1_n10933_25858# vss m1_n10796_25662# vss nfet$221
Xnfet$197_73 m1_13668_17714# vss m1_16538_15778# vss nfet$197
Xnfet$197_62 m1_18665_17343# m1_20721_15778# m1_20104_16080# vss nfet$197
Xnfet$197_51 m1_n7513_20152# vss m1_22493_16080# vss nfet$197
Xpfet$184_1 vdd vdd vdd m1_2822_19850# m1_4620_20152# m1_4620_20152# pfet$184
Xnfet$197_40 m1_n2250_17343# m1_n194_15778# m1_n811_16080# vss nfet$197
Xpfet$206_5 vdd m1_n6839_21786# vdd m1_n5764_21786# pfet$206
Xnfet$212_1 define m1_35837_22102# vss vss nfet$212
Xnfet$205_0 m1_n290_24224# m1_n290_24224# m1_n646_24542# m1_n646_24542# m1_n192_24542#
+ vss nfet$205
Xpfet$181_59 vdd vdd m1_16322_21786# pd6 pfet$181
Xpfet$181_48 vdd m1_16085_25662# m1_15822_23922# m1_15598_25662# pfet$181
Xpfet$181_37 vdd vdd m1_9973_24542# m1_7577_25858# pfet$181
Xpfet$181_26 vdd m1_4997_25658# m1_5790_24542# m1_3049_25662# pfet$181
Xpfet$181_15 vdd m1_11902_25662# m1_11639_23922# m1_11415_25662# pfet$181
Xpfet$211_3 vdd m1_n6839_20152# vdd m1_n927_19404# pfet$211
Xnfet$194_74 pd8 vss m1_23356_21786# vss nfet$194
Xnfet$194_63 m1_14556_21786# vss m1_19644_25858# vss nfet$194
Xnfet$194_52 m1_20126_25858# vss m1_22522_24542# vss nfet$194
Xnfet$194_41 pd5 vss m1_12805_21786# vss nfet$194
Xnfet$194_30 m1_n7513_20152# vss m1_17058_24346# vss nfet$194
Xnfet$213_26 m1_14127_16080# m1_14127_16080# m1_13668_17714# m1_13668_17714# m1_14225_16398#
+ vss nfet$213
Xnfet$213_15 m1_n1989_16202# m1_n1989_16202# vss vss m1_n2507_16398# vss nfet$213
Xpfet$182_91 vdd m1_24287_16080# m1_23820_18030# m1_22848_17343# pfet$182
Xpfet$182_80 vdd vdd m1_15564_15778# m1_15921_16080# pfet$182
Xpfet$187_14 vdd vdd m1_23486_19550# m1_21564_17714# pfet$187
Xnfet$196_7 m1_n7383_17599# m1_n7383_17599# vss vss m1_n63_20470# vss nfet$196
Xnfet$194_4 m1_2912_25858# vss m1_3049_25662# vss nfet$194
Xpfet$193_6 vdd m1_34278_25658# m1_35071_24542# m1_32330_25662# pfet$193
Xpfet$184_26 vdd m1_n1927_20274# m1_n1927_20274# m1_17526_19550# m1_13198_17714# m1_13198_17714#
+ pfet$184
Xpfet$184_15 vdd vdd vdd m1_n59_19550# m1_n7401_15478# m1_n7401_15478# pfet$184
Xpfet$186_5 vdd vdd m1_n6788_16080# m1_n7513_20152# pfet$186
Xnfet$221_6 m1_n10452_25858# vss m1_n10309_25662# vss nfet$221
Xnfet$197_74 m1_14482_17343# vss m1_14641_17836# vss nfet$197
Xnfet$197_63 m1_13668_17714# vss m1_14258_17518# vss nfet$197
Xnfet$197_52 m1_23007_17836# m1_24287_16080# m1_23820_18030# vss nfet$197
Xnfet$207_4 m1_32818_20470# m1_32818_20470# vss vss m1_34329_20470# vss nfet$207
Xnfet$214_5 m1_5148_15478# m1_5148_15478# m1_9624_19404# m1_9624_19404# m1_9856_20470#
+ vss nfet$214
Xnfet$197_30 sd6 vss m1_5148_15478# vss nfet$197
Xnfet$197_41 m1_n2091_17836# m1_n1168_15778# m1_n1989_16202# vss nfet$197
Xpfet$206_6 vdd vdd m1_n6973_21481# m1_n6839_21786# pfet$206
Xpfet$184_2 vdd m1_2590_19404# m1_2590_19404# m1_2822_19850# m1_2384_19550# m1_2384_19550#
+ pfet$184
Xnfet$205_1 m1_814_25658# m1_814_25658# vss vss m1_1273_25502# vss nfet$205
Xpfet$181_49 vdd m1_20126_25858# vdd m1_21729_25658# pfet$181
Xpfet$181_38 vdd vdd m1_16085_25662# m1_15943_25858# pfet$181
Xpfet$181_27 vdd vdd m1_11278_25858# m1_7522_21786# pfet$181
Xpfet$181_16 vdd vdd m1_5771_21786# pd3 pfet$181
Xpfet$211_4 vdd vdd m1_n6839_20152# m1_n6973_21481# pfet$211
Xnfet$194_75 m1_28371_23922# vss m1_28991_24224# vss nfet$194
Xnfet$194_64 m1_19644_25858# vss m1_19781_25662# vss nfet$194
Xnfet$194_53 m1_23827_25858# m1_24451_25662# m1_24188_23922# vss nfet$194
Xnfet$194_42 m1_15943_25858# vss m1_16085_25662# vss nfet$194
Xnfet$194_31 m1_15943_25858# vss m1_18339_24542# vss nfet$194
Xnfet$213_27 m1_18310_16080# m1_18310_16080# vss vss m1_19873_17358# vss nfet$213
Xnfet$213_16 m1_19747_15778# m1_19747_15778# m1_19637_18030# m1_19637_18030# m1_19873_17358#
+ vss nfet$213
Xnfet$194_20 pd3 vss m1_5771_21786# vss nfet$194
Xpfet$182_81 vdd vdd m1_13668_17714# m1_14127_16080# pfet$182
Xpfet$182_70 vdd vdd m1_18824_17836# m1_18665_17343# pfet$182
Xpfet$202_0 vdd vdd vdd m1_n6624_23622# m1_n7082_23622# m1_n7082_23622# pfet$202
Xpfet$182_92 vdd m1_15454_18030# vdd m1_14127_16080# pfet$182
Xpfet$187_15 vdd vdd m1_22205_20152# m1_17697_15478# pfet$187
Xnfet$196_8 m1_27003_19550# m1_27003_19550# vss vss m1_27441_20470# vss nfet$196
Xnfet$194_5 m1_2912_25858# m1_3536_25662# m1_3273_23922# vss nfet$194
Xpfet$193_7 vdd m1_32554_23922# m1_32818_24542# m1_32193_25858# pfet$193
Xpfet$184_27 vdd vdd vdd m1_20407_19850# m1_22205_20152# m1_22205_20152# pfet$184
Xpfet$184_16 vdd vdd vdd m1_28077_19550# m1_26063_15478# m1_26063_15478# pfet$184
Xnfet$228_0 m1_n4485_20152# m1_n6380_21786# vss vss nfet$228
Xpfet$186_6 vdd vdd m1_n7383_17599# m1_n7247_17714# pfet$186
Xpfet$207_10 vdd vdd m1_n10933_25858# fin pfet$207
Xnfet$197_75 sd3 vss m1_17697_15478# vss nfet$197
Xnfet$197_64 m1_13668_17714# vss m1_13198_17714# vss nfet$197
Xnfet$197_53 m1_22848_17343# vss m1_23007_17836# vss nfet$197
Xnfet$207_5 m1_32818_21586# m1_32818_21586# m1_34093_19792# m1_34093_19792# m1_34329_20470#
+ vss nfet$207
Xnfet$197_31 m1_1933_17343# m1_3989_15778# m1_3372_16080# vss nfet$197
Xnfet$197_20 m1_1119_17714# vss m1_1709_17518# vss nfet$197
Xnfet$214_6 m1_11654_20152# m1_11654_20152# m1_9624_19404# m1_9624_19404# m1_10488_20470#
+ vss nfet$214
Xnfet$197_42 m1_n811_16080# vss m1_n1168_15778# vss nfet$197
Xnfet$221_7 m1_n7320_25516# vss m1_n2567_23922# vss nfet$221
Xpfet$206_7 vdd vdd m1_n6839_21786# m1_n6380_21786# pfet$206
Xpfet$184_3 vdd vdd vdd m1_3458_19550# m1_n3218_15478# m1_n3218_15478# pfet$184
Xnfet$205_2 m1_326_24346# m1_326_24346# m1_n789_25858# m1_n789_25858# m1_1273_25502#
+ vss nfet$205
Xpfet$181_39 vdd vdd m1_15598_25662# m1_15461_25858# pfet$181
Xpfet$181_28 vdd m1_11639_23922# m1_11903_24542# m1_11278_25858# pfet$181
Xpfet$181_17 vdd vdd m1_7577_25858# m1_8692_24346# pfet$181
Xpfet$182_0 vdd vdd m1_12355_15778# m1_9485_17714# pfet$182
Xnfet$194_76 m1_28492_25858# vss m1_28634_25662# vss nfet$194
Xnfet$194_65 m1_28492_25858# vss m1_25107_21786# vss nfet$194
Xnfet$194_54 m1_24309_25858# vss m1_24451_25662# vss nfet$194
Xnfet$194_43 m1_15461_25858# vss m1_15598_25662# vss nfet$194
Xnfet$194_32 m1_15461_25858# m1_17546_25658# m1_18339_24542# vss nfet$194
Xnfet$213_17 m1_22493_16080# m1_22493_16080# vss vss m1_24056_17358# vss nfet$213
Xnfet$210_0 m1_34093_19792# vss m1_34843_21786# vss nfet$210
Xnfet$194_21 m1_11278_25858# m1_11902_25662# m1_11639_23922# vss nfet$194
Xnfet$194_10 m1_7577_25858# vss m1_9973_24542# vss nfet$194
Xpfet$202_1 vdd m1_n6856_24542# m1_n6856_24542# m1_n6624_23622# m1_n8283_19850# m1_n8283_19850#
+ pfet$202
Xpfet$182_93 vdd m1_23820_18030# vdd m1_22493_16080# pfet$182
Xpfet$182_82 vdd m1_13668_17714# vdd m1_14743_16202# pfet$182
Xpfet$182_71 vdd vdd m1_19747_15778# m1_20104_16080# pfet$182
Xpfet$182_60 vdd vdd m1_n194_15778# m1_n3064_17714# pfet$182
Xpfet$187_16 vdd vdd m1_19969_19550# m1_17381_17714# pfet$187
Xnfet$196_9 m1_25747_17714# m1_25747_17714# vss vss m1_28073_20470# vss nfet$196
Xpfet$186_7 vdd vdd m1_27190_17836# m1_27031_17343# pfet$186
Xnfet$194_6 m1_3049_25662# m1_3893_24224# m1_4997_25658# vss nfet$194
Xnfet$228_1 m1_n5227_20152# vss m1_n6380_21786# vss nfet$228
Xpfet$207_11 vdd vdd m1_n9336_24346# vss pfet$207
Xpfet$184_28 vdd vdd vdd m1_21043_19550# m1_17697_15478# m1_17697_15478# pfet$184
Xpfet$184_17 vdd m1_n3822_20130# m1_n3822_20130# m1_28077_19550# m1_25747_17714# m1_25747_17714#
+ pfet$184
Xnfet$207_6 m1_354_22513# m1_354_22513# m1_31535_22102# m1_31535_22102# m1_31771_21430#
+ vss nfet$207
Xnfet$214_7 m1_n7401_15478# m1_n7401_15478# m1_n927_19404# m1_n927_19404# m1_n695_20470#
+ vss nfet$214
Xnfet$197_10 m1_11738_16080# vss m1_11381_15778# vss nfet$197
Xnfet$221_8 m1_n4623_25487# vss m1_n4464_25980# vss nfet$221
Xnfet$197_76 m1_14482_17343# m1_16538_15778# m1_15921_16080# vss nfet$197
Xnfet$197_65 m1_14482_17343# m1_14743_16202# m1_14258_17518# vss nfet$197
Xnfet$197_54 m1_22848_17343# m1_23109_16202# m1_22624_17518# vss nfet$197
Xpfet$184_4 vdd m1_6107_19404# m1_6107_19404# m1_6339_19850# m1_5901_19550# m1_5901_19550#
+ pfet$184
Xnfet$197_32 m1_2092_17836# m1_3015_15778# m1_2194_16202# vss nfet$197
Xnfet$197_21 m1_1933_17343# m1_2194_16202# m1_1709_17518# vss nfet$197
Xnfet$197_43 sd8 vss m1_n3218_15478# vss nfet$197
Xnfet$205_3 m1_326_24346# m1_326_24346# vss vss m1_n192_24542# vss nfet$205
Xpfet$181_29 vdd vdd m1_11903_24542# m1_12259_24224# pfet$181
Xpfet$181_18 vdd vdd m1_11415_25662# m1_11278_25858# pfet$181
Xpfet$182_1 vdd vdd m1_11381_15778# m1_11738_16080# pfet$182
Xnfet$194_77 m1_28010_25858# vss m1_28147_25662# vss nfet$194
Xnfet$194_66 m1_28010_25858# m1_30095_25658# m1_30888_24542# vss nfet$194
Xnfet$194_55 m1_23827_25858# vss m1_23964_25662# vss nfet$194
Xnfet$194_44 m1_15822_23922# vss m1_16442_24224# vss nfet$194
Xnfet$194_33 m1_11760_25858# vss m1_14156_24542# vss nfet$194
Xnfet$210_1 m1_30256_19792# vss m1_32818_20470# vss nfet$210
Xnfet$194_22 m1_11760_25858# vss m1_11902_25662# vss nfet$194
Xnfet$194_11 m1_7522_21786# vss m1_11278_25858# vss nfet$194
Xnfet$203_0 m1_n1134_25662# m1_n910_23922# m1_n646_24542# vss nfet$203
Xnfet$213_18 m1_23930_15778# m1_23930_15778# m1_23820_18030# m1_23820_18030# m1_24056_17358#
+ vss nfet$213
Xpfet$182_94 vdd vdd m1_22624_17518# m1_22034_17714# pfet$182
Xpfet$182_83 vdd m1_16538_15778# m1_15921_16080# m1_14641_17836# pfet$182
Xpfet$182_72 vdd m1_20721_15778# m1_20104_16080# m1_18824_17836# pfet$182
Xpfet$182_61 vdd m1_n811_16080# m1_n1278_18030# m1_n2250_17343# pfet$182
Xpfet$182_50 vdd m1_n1168_15778# m1_n1989_16202# m1_n2250_17343# pfet$182
Xpfet$187_17 vdd vdd m1_25722_20152# m1_21880_15478# pfet$187
Xnfet$194_7 m1_3049_25662# m1_3273_23922# m1_3537_24542# vss nfet$194
Xpfet$207_12 vdd vdd m1_n7082_23622# m1_n8625_26174# pfet$207
Xpfet$184_29 vdd vdd vdd m1_23924_19850# m1_25722_20152# m1_25722_20152# pfet$184
Xpfet$184_18 vdd vdd vdd m1_27441_19850# m1_29239_20152# m1_29239_20152# pfet$184
Xpfet$186_8 vdd vdd m1_28113_15778# m1_28470_16080# pfet$186
Xnfet$207_7 m1_3871_22513# m1_3871_22513# vss vss m1_31771_21430# vss nfet$207
Xnfet$214_8 m1_26063_15478# m1_26063_15478# m1_n3822_20130# m1_n3822_20130# m1_27441_20470#
+ vss nfet$214
Xnfet$221_9 m1_n3184_24224# vss m1_n3541_23922# vss nfet$221
Xnfet$197_77 sd4 vss m1_13514_15478# vss nfet$197
Xnfet$197_66 m1_n7513_20152# vss m1_14127_16080# vss nfet$197
Xnfet$197_55 m1_22034_17714# vss m1_24904_15778# vss nfet$197
Xnfet$197_44 m1_n2091_17836# m1_n811_16080# m1_n1278_18030# vss nfet$197
Xpfet$184_5 vdd vdd vdd m1_n695_19850# m1_1103_20152# m1_1103_20152# pfet$184
Xnfet$197_33 sd7 vss m1_965_15478# vss nfet$197
Xnfet$197_22 m1_6116_17343# m1_6377_16202# m1_5892_17518# vss nfet$197
Xnfet$197_11 m1_10299_17343# m1_12355_15778# m1_11738_16080# vss nfet$197
Xnfet$205_4 m1_33174_24224# m1_33174_24224# m1_32818_24542# m1_32818_24542# m1_33272_24542#
+ vss nfet$205
Xpfet$181_19 vdd vdd m1_7095_25858# m1_4005_21786# pfet$181
Xpfet$182_2 vdd m1_12355_15778# m1_11738_16080# m1_10458_17836# pfet$182
Xnfet$194_78 m1_28010_25858# m1_28634_25662# m1_28371_23922# vss nfet$194
Xnfet$194_67 m1_28492_25858# vss m1_30888_24542# vss nfet$194
Xnfet$194_56 m1_19781_25662# m1_20625_24224# m1_21729_25658# vss nfet$194
Xnfet$194_45 m1_15461_25858# m1_16085_25662# m1_15822_23922# vss nfet$194
Xnfet$194_34 m1_11278_25858# m1_13363_25658# m1_14156_24542# vss nfet$194
Xnfet$210_2 m1_31535_19792# m1_32818_20470# vss vss nfet$210
Xnfet$194_23 m1_11278_25858# vss m1_11415_25662# vss nfet$194
Xnfet$194_12 m1_7577_25858# vss m1_7522_21786# vss nfet$194
Xnfet$213_19 m1_23109_16202# m1_23109_16202# vss vss m1_22591_16398# vss nfet$213
Xnfet$203_1 m1_n1271_25858# m1_n647_25662# m1_n910_23922# vss nfet$203
Xpfet$182_95 vdd vdd m1_21564_17714# m1_22034_17714# pfet$182
Xpfet$182_84 vdd vdd m1_17381_17714# m1_17851_17714# pfet$182
Xpfet$182_73 vdd vdd m1_16538_15778# m1_13668_17714# pfet$182
Xpfet$182_62 vdd vdd m1_23007_17836# m1_22848_17343# pfet$182
Xpfet$182_40 vdd m1_10560_16202# m1_10075_17518# m1_10458_17836# pfet$182
Xpfet$182_51 vdd vdd m1_n1168_15778# m1_n811_16080# pfet$182
Xpfet$200_0 vdd m1_n4377_15778# m1_n4994_16080# m1_n6274_17836# pfet$200
Xnfet$194_8 m1_3394_25858# vss m1_3536_25662# vss nfet$194
Xpfet$207_13 vdd vdd m1_n8055_24542# m1_n8625_26174# pfet$207
Xpfet$184_19 vdd m1_n3822_20130# m1_n3822_20130# m1_27441_19850# m1_27003_19550# m1_27003_19550#
+ pfet$184
Xpfet$186_9 vdd vdd m1_29087_15778# m1_26217_17714# pfet$186
Xpfet$198_0 vdd m1_32818_20470# m1_32818_20470# m1_33050_19550# m1_30256_19792# m1_30256_19792#
+ pfet$198
Xnfet$214_9 m1_29239_20152# m1_29239_20152# m1_n3822_20130# m1_n3822_20130# m1_28073_20470#
+ vss nfet$214
Xnfet$197_78 m1_14641_17836# m1_15564_15778# m1_14743_16202# vss nfet$197
Xnfet$197_67 m1_17381_17714# vss m1_14482_17343# vss nfet$197
Xnfet$197_56 m1_24287_16080# vss m1_23930_15778# vss nfet$197
Xnfet$197_45 m1_n3064_17714# vss m1_n194_15778# vss nfet$197
Xnfet$197_34 m1_n2250_17343# vss m1_n2091_17836# vss nfet$197
Xnfet$197_23 m1_5302_17714# vss m1_4832_17714# vss nfet$197
Xnfet$197_12 m1_9485_17714# vss m1_12355_15778# vss nfet$197
Xpfet$184_6 vdd vdd vdd m1_6339_19850# m1_8137_20152# m1_8137_20152# pfet$184
Xnfet$226_0 m1_n4485_21904# m1_n5764_21786# vss vss nfet$226
Xnfet$205_5 m1_33790_24346# m1_33790_24346# vss vss m1_33272_24542# vss nfet$205
Xpfet$182_3 vdd m1_11381_15778# m1_10560_16202# m1_10299_17343# pfet$182
Xnfet$194_79 pd7 vss m1_19839_21786# vss nfet$194
Xnfet$194_68 m1_n7513_20152# vss m1_29607_24346# vss nfet$194
Xnfet$210_3 m1_30256_22102# vss m1_32818_21586# vss nfet$210
Xnfet$194_57 m1_20126_25858# vss m1_20268_25662# vss nfet$194
Xnfet$194_46 m1_20126_25858# vss m1_18073_21786# vss nfet$194
Xnfet$194_35 m1_15598_25662# m1_15822_23922# m1_16086_24542# vss nfet$194
Xnfet$194_24 m1_7095_25858# m1_7719_25662# m1_7456_23922# vss nfet$194
Xnfet$194_13 m1_11415_25662# m1_11639_23922# m1_11903_24542# vss nfet$194
Xnfet$203_2 m1_n1271_25858# m1_814_25658# m1_1607_24542# vss nfet$203
Xpfet$182_96 vdd vdd m1_18665_17343# m1_21564_17714# pfet$182
Xpfet$182_85 vdd m1_18926_16202# m1_18441_17518# m1_18824_17836# pfet$182
Xpfet$182_74 vdd vdd m1_14641_17836# m1_14482_17343# pfet$182
Xpfet$182_63 vdd m1_23930_15778# m1_23109_16202# m1_22848_17343# pfet$182
Xpfet$182_30 vdd vdd m1_1933_17343# m1_4832_17714# pfet$182
Xpfet$182_41 vdd vdd m1_10075_17518# m1_9485_17714# pfet$182
Xpfet$182_52 vdd m1_n3064_17714# vdd m1_n1989_16202# pfet$182
Xpfet$200_1 vdd m1_n5351_15778# m1_n6172_16202# m1_n6433_17343# pfet$200
Xnfet$194_9 m1_3273_23922# vss m1_3893_24224# vss nfet$194
Xpfet$198_1 vdd vdd vdd m1_33050_19550# m1_31535_19792# m1_31535_19792# pfet$198
Xnfet$197_79 m1_15921_16080# vss m1_15564_15778# vss nfet$197
Xnfet$197_68 m1_18665_17343# m1_18926_16202# m1_18441_17518# vss nfet$197
Xnfet$197_57 m1_22848_17343# m1_24904_15778# m1_24287_16080# vss nfet$197
Xnfet$197_46 m1_22034_17714# vss m1_21564_17714# vss nfet$197
Xnfet$197_24 m1_4832_17714# vss m1_1933_17343# vss nfet$197
Xnfet$197_13 m1_10458_17836# m1_11381_15778# m1_10560_16202# vss nfet$197
Xnfet$197_35 m1_n7513_20152# vss m1_5761_16080# vss nfet$197
Xnfet$226_1 m1_n5227_21418# vss m1_n5764_21786# vss nfet$226
Xnfet$219_0 m1_n7082_23622# m1_n6856_24542# vss vss nfet$219
Xpfet$182_110 vdd vdd m1_10458_17836# m1_10299_17343# pfet$182
Xpfet$184_7 vdd vdd vdd m1_6975_19550# m1_965_15478# m1_965_15478# pfet$184
Xnfet$205_6 m1_33790_24346# m1_33790_24346# m1_32675_25947# m1_32675_25947# m1_34737_25502#
+ vss nfet$205
Xpfet$182_4 vdd m1_9485_17714# vdd m1_10560_16202# pfet$182
Xnfet$194_69 m1_24309_25858# vss m1_26705_24542# vss nfet$194
Xnfet$194_58 m1_20005_23922# vss m1_20625_24224# vss nfet$194
Xnfet$194_47 m1_23964_25662# m1_24188_23922# m1_24452_24542# vss nfet$194
Xnfet$194_36 m1_11760_25858# vss m1_11039_21786# vss nfet$194
Xnfet$194_25 m1_7232_25662# m1_8076_24224# m1_9180_25658# vss nfet$194
Xnfet$194_14 m1_n7513_20152# vss m1_8692_24346# vss nfet$194
Xnfet$203_3 m1_n1134_25662# m1_n290_24224# m1_814_25658# vss nfet$203
Xpfet$182_97 vdd vdd m1_22493_16080# m1_n7513_20152# pfet$182
Xpfet$182_86 vdd m1_19637_18030# vdd m1_18310_16080# pfet$182
Xpfet$182_75 vdd vdd m1_17697_15478# sd3 pfet$182
Xpfet$182_64 vdd vdd m1_23930_15778# m1_24287_16080# pfet$182
Xpfet$182_20 vdd vdd m1_1119_17714# m1_1578_16080# pfet$182
Xpfet$182_31 vdd m1_3372_16080# m1_2905_18030# m1_1933_17343# pfet$182
Xpfet$182_42 vdd m1_11271_18030# vdd m1_9944_16080# pfet$182
Xpfet$182_53 vdd vdd m1_n3218_15478# sd8 pfet$182
Xnfet$201_0 m1_n3534_17714# vss m1_n6433_17343# vss nfet$201
Xpfet$200_2 vdd m1_n4994_16080# m1_n5461_18030# m1_n6433_17343# pfet$200
Xnfet$199_0 m1_n3534_17714# vss m1_2384_19550# vss nfet$199
Xpfet$198_2 vdd m1_32818_21586# m1_32818_21586# m1_33050_22344# m1_30256_22102# m1_30256_22102#
+ pfet$198
Xnfet$197_69 m1_17851_17714# vss m1_17381_17714# vss nfet$197
Xnfet$197_58 m1_23007_17836# m1_23930_15778# m1_23109_16202# vss nfet$197
Xnfet$197_47 m1_22034_17714# vss m1_22624_17518# vss nfet$197
Xnfet$197_25 m1_2092_17836# m1_3372_16080# m1_2905_18030# vss nfet$197
Xnfet$197_14 m1_6116_17343# m1_8172_15778# m1_7555_16080# vss nfet$197
Xnfet$197_36 m1_n3064_17714# vss m1_n2474_17518# vss nfet$197
Xpfet$184_8 vdd m1_9624_19404# m1_9624_19404# m1_10492_19550# m1_4832_17714# m1_4832_17714#
+ pfet$184
Xnfet$226_2 m1_n6839_21786# vss m1_n6973_21481# vss nfet$226
Xnfet$219_1 m1_n8283_19850# vss m1_n6856_24542# vss nfet$219
Xnfet$205_7 m1_34278_25658# m1_34278_25658# vss vss m1_34737_25502# vss nfet$205
Xnfet$206_10 m1_21590_21786# m1_21590_21786# vss vss m1_20428_21586# vss nfet$206
Xpfet$182_100 vdd vdd m1_23820_18030# m1_23930_15778# pfet$182
Xpfet$182_5 vdd m1_7198_15778# m1_6377_16202# m1_6116_17343# pfet$182
Xnfet$203_4 m1_32193_25858# m1_34278_25658# m1_35071_24542# vss nfet$203
Xnfet$194_59 m1_19644_25858# m1_20268_25662# m1_20005_23922# vss nfet$194
Xnfet$194_48 m1_18073_21786# vss m1_23827_25858# vss nfet$194
Xnfet$194_37 m1_11039_21786# vss m1_15461_25858# vss nfet$194
Xnfet$194_26 m1_7095_25858# m1_9180_25658# m1_9973_24542# vss nfet$194
Xnfet$194_15 m1_7232_25662# m1_7456_23922# m1_7720_24542# vss nfet$194
Xpfet$182_98 vdd m1_20104_16080# m1_19637_18030# m1_18665_17343# pfet$182
Xpfet$182_87 vdd vdd m1_18310_16080# m1_n7513_20152# pfet$182
Xpfet$182_76 vdd m1_17851_17714# vdd m1_18926_16202# pfet$182
Xpfet$182_65 vdd m1_24904_15778# m1_24287_16080# m1_23007_17836# pfet$182
Xpfet$182_21 vdd vdd m1_965_15478# sd7 pfet$182
Xpfet$182_10 vdd m1_8172_15778# m1_7555_16080# m1_6275_17836# pfet$182
Xpfet$182_32 vdd vdd m1_2905_18030# m1_3015_15778# pfet$182
Xpfet$182_43 vdd vdd m1_11271_18030# m1_11381_15778# pfet$182
Xpfet$182_54 vdd vdd m1_n1278_18030# m1_n1168_15778# pfet$182
Xnfet$201_1 m1_n7513_20152# vss m1_n6788_16080# vss nfet$201
Xpfet$200_3 vdd m1_n6172_16202# m1_n6657_17518# m1_n6274_17836# pfet$200
Xnfet$214_10 m1_9331_15478# m1_9331_15478# m1_n3822_21786# m1_n3822_21786# m1_13373_20470#
+ vss nfet$214
Xnfet$199_1 m1_n3218_15478# vss m1_4620_20152# vss nfet$199
Xnfet$197_15 m1_5302_17714# vss m1_8172_15778# vss nfet$197
Xnfet$197_59 m1_17851_17714# vss m1_20721_15778# vss nfet$197
Xnfet$197_48 m1_18824_17836# m1_20104_16080# m1_19637_18030# vss nfet$197
Xnfet$197_26 m1_5302_17714# vss m1_5892_17518# vss nfet$197
Xpfet$184_9 vdd m1_9624_19404# m1_9624_19404# m1_9856_19850# m1_9418_19550# m1_9418_19550#
+ pfet$184
Xnfet$197_37 m1_n7513_20152# vss m1_n2605_16080# vss nfet$197
Xpfet$196_0 vdd vdd vdd m1_36073_22344# define define pfet$196
Xpfet$185_10 vdd vdd m1_23486_21590# m1_23356_21786# pfet$185
Xnfet$206_11 m1_22222_21786# m1_22222_21786# vss vss m1_21060_21586# vss nfet$206
Xpfet$182_101 vdd vdd m1_19637_18030# m1_19747_15778# pfet$182
Xnfet$224_0 m1_n7186_25858# vss m1_n7320_25516# vss nfet$224
Xpfet$182_6 vdd vdd m1_7198_15778# m1_7555_16080# pfet$182
Xpfet$209_0 vdd vdd vdd m1_n8047_19550# m1_n7513_20152# m1_n7513_20152# pfet$209
Xnfet$203_5 m1_32330_25662# m1_33174_24224# m1_34278_25658# vss nfet$203
Xnfet$194_49 m1_19781_25662# m1_20005_23922# m1_20269_24542# vss nfet$194
Xnfet$194_38 m1_n7513_20152# vss m1_12875_24346# vss nfet$194
Xnfet$194_27 m1_7577_25858# vss m1_7719_25662# vss nfet$194
Xnfet$194_16 m1_4005_21786# vss m1_7095_25858# vss nfet$194
Xpfet$182_99 vdd m1_23109_16202# m1_22624_17518# m1_23007_17836# pfet$182
Xpfet$182_88 vdd vdd m1_18441_17518# m1_17851_17714# pfet$182
Xpfet$182_77 vdd vdd m1_17851_17714# m1_18310_16080# pfet$182
Xpfet$182_66 vdd vdd m1_24904_15778# m1_22034_17714# pfet$182
Xpfet$182_22 vdd vdd m1_3015_15778# m1_3372_16080# pfet$182
Xpfet$182_11 vdd vdd m1_9485_17714# m1_9944_16080# pfet$182
Xpfet$182_33 vdd vdd m1_5892_17518# m1_5302_17714# pfet$182
Xpfet$182_44 vdd vdd m1_649_17714# m1_1119_17714# pfet$182
Xpfet$182_55 vdd vdd m1_n2474_17518# m1_n3064_17714# pfet$182
Xnfet$201_2 m1_n4994_16080# vss m1_n5351_15778# vss nfet$201
Xnfet$214_11 m1_15171_20152# m1_15171_20152# m1_n3822_21786# m1_n3822_21786# m1_14005_20470#
+ vss nfet$214
Xpfet$200_4 vdd m1_28113_15778# m1_27292_16202# m1_27031_17343# pfet$200
Xnfet$199_2 m1_n7401_15478# vss m1_1103_20152# vss nfet$199
Xnfet$197_49 m1_21564_17714# vss m1_18665_17343# vss nfet$197
Xnfet$197_27 m1_1119_17714# vss m1_3989_15778# vss nfet$197
Xnfet$197_16 m1_6275_17836# m1_7198_15778# m1_6377_16202# vss nfet$197
Xnfet$197_38 m1_n2250_17343# m1_n1989_16202# m1_n2474_17518# vss nfet$197
Xpfet$196_1 vdd m1_35837_22102# m1_35837_22102# m1_36073_22344# fout fout pfet$196
Xpfet$185_11 vdd vdd m1_18705_21786# m1_18073_21786# pfet$185
Xnfet$206_12 m1_18073_21786# m1_18073_21786# vss vss m1_16911_21586# vss nfet$206
Xpfet$182_102 vdd vdd m1_13198_17714# m1_13668_17714# pfet$182
Xpfet$189_0 vdd vdd m1_n647_25662# m1_n789_25858# pfet$189
Xpfet$182_7 vdd vdd m1_6275_17836# m1_6116_17343# pfet$182
Xnfet$217_0 m1_n5351_15778# m1_n5351_15778# m1_n5461_18030# m1_n5461_18030# m1_n5225_17358#
+ vss nfet$217
Xpfet$209_1 vdd m1_n8283_19850# m1_n8283_19850# m1_n8047_19550# m1_n8283_20611# m1_n8283_20611#
+ pfet$209
Xnfet$224_1 m1_n6856_24542# vss m1_n6111_25858# vss nfet$224
Xnfet$194_39 pd4 vss m1_9288_21786# vss nfet$194
Xnfet$194_28 m1_3394_25858# vss m1_4005_21786# vss nfet$194
Xnfet$194_17 m1_11639_23922# vss m1_12259_24224# vss nfet$194
Xnfet$203_6 m1_32193_25858# m1_32817_25662# m1_32554_23922# vss nfet$203
Xpfet$182_89 vdd vdd m1_22848_17343# m1_25747_17714# pfet$182
Xpfet$182_78 vdd vdd m1_13514_15478# sd4 pfet$182
Xpfet$182_67 vdd m1_22034_17714# vdd m1_23109_16202# pfet$182
Xpfet$182_12 vdd m1_3989_15778# m1_3372_16080# m1_2092_17836# pfet$182
Xpfet$182_23 vdd m1_5302_17714# vdd m1_6377_16202# pfet$182
Xpfet$182_34 vdd vdd m1_5761_16080# m1_n7513_20152# pfet$182
Xpfet$182_45 vdd vdd m1_9944_16080# m1_n7513_20152# pfet$182
Xpfet$182_56 vdd m1_n1278_18030# vdd m1_n2605_16080# pfet$182
Xnfet$201_3 m1_n6433_17343# vss m1_n6274_17836# vss nfet$201
Xnfet$214_12 m1_18688_20152# m1_18688_20152# m1_n1927_20274# m1_n1927_20274# m1_17522_20470#
+ vss nfet$214
Xpfet$200_5 vdd m1_29087_15778# m1_28470_16080# m1_27190_17836# pfet$200
Xnfet$199_3 m1_649_17714# vss m1_5901_19550# vss nfet$199
Xnfet$197_28 m1_1933_17343# vss m1_2092_17836# vss nfet$197
Xnfet$197_17 m1_649_17714# vss m1_n2250_17343# vss nfet$197
Xnfet$197_39 m1_n3064_17714# vss m1_n3534_17714# vss nfet$197
Xpfet$185_12 vdd vdd m1_16452_21590# m1_16322_21786# pfet$185
Xnfet$206_13 m1_18705_21786# m1_18705_21786# vss vss m1_17543_21586# vss nfet$206
Xpfet$182_103 vdd m1_14743_16202# m1_14258_17518# m1_14641_17836# pfet$182
Xnfet$197_0 m1_9485_17714# vss m1_9015_17714# vss nfet$197
Xpfet$189_1 vdd vdd m1_n1134_25662# m1_n1271_25858# pfet$189
Xpfet$182_8 vdd vdd m1_9331_15478# sd5 pfet$182
Xnfet$217_1 m1_n6788_16080# m1_n6788_16080# vss vss m1_n5225_17358# vss nfet$217
Xpfet$209_2 vdd m1_n8283_20611# m1_n8283_20611# m1_n8047_22344# m1_n8145_21908# m1_n8145_21908#
+ pfet$209
Xnfet$203_7 m1_32330_25662# m1_32554_23922# m1_32818_24542# vss nfet$203
Xnfet$194_29 m1_15943_25858# vss m1_14556_21786# vss nfet$194
Xnfet$194_18 m1_7095_25858# vss m1_7232_25662# vss nfet$194
Xpfet$182_79 vdd m1_15564_15778# m1_14743_16202# m1_14482_17343# pfet$182
Xpfet$182_68 vdd vdd m1_22034_17714# m1_22493_16080# pfet$182
Xpfet$182_13 vdd vdd m1_5148_15478# sd6 pfet$182
Xpfet$182_24 vdd m1_6377_16202# m1_5892_17518# m1_6275_17836# pfet$182
Xpfet$182_35 vdd vdd m1_9015_17714# m1_9485_17714# pfet$182
Xpfet$182_46 vdd vdd m1_n2250_17343# m1_649_17714# pfet$182
Xpfet$182_57 vdd m1_n1989_16202# m1_n2474_17518# m1_n2091_17836# pfet$182
Xnfet$201_4 m1_n7247_17714# vss m1_n4377_15778# vss nfet$201
Xnfet$214_13 m1_13514_15478# m1_13514_15478# m1_n1927_20274# m1_n1927_20274# m1_16890_20470#
+ vss nfet$214
Xpfet$200_6 vdd m1_28470_16080# m1_28003_18030# m1_27031_17343# pfet$200
Xnfet$199_4 m1_4832_17714# vss m1_9418_19550# vss nfet$199
Xnfet$197_29 m1_3372_16080# vss m1_3015_15778# vss nfet$197
Xnfet$197_18 m1_1119_17714# vss m1_649_17714# vss nfet$197
Xnfet$206_14 m1_15188_21786# m1_15188_21786# vss vss m1_14026_21586# vss nfet$206
Xpfet$182_104 vdd vdd m1_14127_16080# m1_n7513_20152# pfet$182
Xnfet$197_1 m1_9015_17714# vss m1_6116_17343# vss nfet$197
Xpfet$189_2 vdd vdd m1_n1271_25858# m1_n10452_25858# pfet$189
Xpfet$185_13 vdd vdd m1_15188_21786# m1_14556_21786# pfet$185
Xpfet$182_9 vdd vdd m1_8172_15778# m1_5302_17714# pfet$182
Xnfet$217_2 m1_n6788_16080# m1_n6788_16080# m1_n7247_17714# m1_n7247_17714# m1_n6690_16398#
+ vss nfet$217
Xpfet$194_0 vdd vdd m1_n1263_21786# pd1 pfet$194
Xpfet$209_3 vdd vdd vdd m1_n8047_22344# m1_n8283_19850# m1_n8283_19850# pfet$209
Xnfet$194_19 m1_7456_23922# vss m1_8076_24224# vss nfet$194
Xpfet$182_69 vdd vdd m1_20721_15778# m1_17851_17714# pfet$182
Xpfet$182_14 vdd vdd m1_2092_17836# m1_1933_17343# pfet$182
Xpfet$182_25 vdd vdd m1_1709_17518# m1_1119_17714# pfet$182
Xpfet$182_36 vdd vdd m1_6116_17343# m1_9015_17714# pfet$182
Xpfet$182_47 vdd m1_11738_16080# m1_11271_18030# m1_10299_17343# pfet$182
Xpfet$182_58 vdd vdd m1_n3534_17714# m1_n3064_17714# pfet$182
Xnfet$222_0 m1_n9952_24224# m1_n9952_24224# m1_n10308_24542# m1_n10308_24542# m1_n9854_24542#
+ vss nfet$222
Xpfet$207_0 vdd vdd m1_n10796_25662# m1_n10933_25858# pfet$207
Xpfet$200_7 vdd m1_27292_16202# m1_26807_17518# m1_27190_17836# pfet$200
Xnfet$201_5 m1_n7247_17714# vss m1_n6657_17518# vss nfet$201
Xnfet$214_14 m1_22205_20152# m1_22205_20152# m1_n2543_20130# m1_n2543_20130# m1_21039_20470#
+ vss nfet$214
Xnfet$199_5 m1_965_15478# vss m1_8137_20152# vss nfet$199
Xnfet$197_19 m1_n7513_20152# vss m1_1578_16080# vss nfet$197
Xnfet$197_2 m1_6275_17836# m1_7555_16080# m1_7088_18030# vss nfet$197
Xpfet$185_14 vdd vdd m1_19969_21590# m1_19839_21786# pfet$185
Xnfet$206_15 m1_14556_21786# m1_14556_21786# vss vss m1_13394_21586# vss nfet$206
Xpfet$182_105 vdd vdd m1_14258_17518# m1_13668_17714# pfet$182
Xpfet$189_3 vdd vdd m1_1607_24542# m1_n789_25858# pfet$189
Xnfet$217_3 m1_n6172_16202# m1_n6172_16202# vss vss m1_n6690_16398# vss nfet$217
Xpfet$194_1 vdd vdd m1_2254_21786# pd2 pfet$194
Xpfet$187_0 vdd vdd m1_2384_19550# m1_n3534_17714# pfet$187
Xnfet$215_0 m1_35837_22102# vss m1_n7513_20152# vss nfet$215
Xnfet$222_1 m1_n9336_24346# m1_n9336_24346# m1_n8625_26174# m1_n8625_26174# m1_n8389_25502#
+ vss nfet$222
Xpfet$182_15 vdd vdd m1_5302_17714# m1_5761_16080# pfet$182
Xpfet$182_26 vdd vdd m1_4832_17714# m1_5302_17714# pfet$182
Xpfet$182_37 vdd m1_7555_16080# m1_7088_18030# m1_6116_17343# pfet$182
Xpfet$182_48 vdd vdd m1_n3064_17714# m1_n2605_16080# pfet$182
Xpfet$182_59 vdd vdd m1_n2605_16080# m1_n7513_20152# pfet$182
Xpfet$207_1 vdd vdd m1_n10309_25662# m1_n10452_25858# pfet$207
Xnfet$201_6 m1_n7247_17714# vss m1_n7383_17599# vss nfet$201
Xnfet$214_15 m1_17697_15478# m1_17697_15478# m1_n2543_20130# m1_n2543_20130# m1_20407_20470#
+ vss nfet$214
Xnfet$199_6 m1_9015_17714# vss m1_12935_19550# vss nfet$199
Xnfet$197_3 m1_n7513_20152# vss m1_9944_16080# vss nfet$197
Xpfet$185_15 vdd vdd m1_27003_21590# m1_26873_21786# pfet$185
Xnfet$206_16 m1_28624_21786# m1_28624_21786# vss vss m1_27462_21586# vss nfet$206
Xpfet$182_106 vdd vdd m1_14482_17343# m1_17381_17714# pfet$182
Xpfet$189_4 vdd vdd m1_488_21786# m1_n789_25858# pfet$189
Xnfet$217_4 m1_28113_15778# m1_28113_15778# m1_28003_18030# m1_28003_18030# m1_28239_17358#
+ vss nfet$217
Xpfet$194_2 vdd vdd m1_26873_21786# pd9 pfet$194
Xnfet$195_0 m1_n1133_21590# m1_n1133_21590# m1_354_22513# m1_354_22513# m1_n674_21586#
+ vss nfet$195
Xpfet$187_1 vdd vdd m1_4620_20152# m1_n3218_15478# pfet$187
Xnfet$208_0 m1_34843_21786# m1_34843_21786# m1_34093_22102# m1_34093_22102# m1_34329_21430#
+ vss nfet$208
Xnfet$222_2 m1_n8848_25658# m1_n8848_25658# vss vss m1_n8389_25502# vss nfet$222
Xpfet$182_16 vdd vdd m1_3989_15778# m1_1119_17714# pfet$182
Xpfet$182_27 vdd m1_2194_16202# m1_1709_17518# m1_2092_17836# pfet$182
Xpfet$182_38 vdd vdd m1_7088_18030# m1_7198_15778# pfet$182
Xpfet$182_49 vdd m1_n194_15778# m1_n811_16080# m1_n2091_17836# pfet$182
Xpfet$207_2 vdd vdd m1_n9952_24224# m1_n10572_23922# pfet$207
Xnfet$201_7 m1_26217_17714# vss m1_26807_17518# vss nfet$201
Xnfet$214_16 m1_25722_20152# m1_25722_20152# m1_n3206_20274# m1_n3206_20274# m1_24556_20470#
+ vss nfet$214
Xpfet$212_0 vdd vdd vdd m1_n5019_19550# m1_n4485_20152# m1_n4485_20152# pfet$212
Xnfet$199_7 m1_5148_15478# vss m1_11654_20152# vss nfet$199
Xnfet$197_4 m1_10299_17343# m1_10560_16202# m1_10075_17518# vss nfet$197
Xpfet$185_16 vdd vdd m1_29256_21786# m1_28624_21786# pfet$185
Xnfet$206_17 m1_29256_21786# m1_29256_21786# vss vss m1_28094_21586# vss nfet$206
Xpfet$182_107 vdd m1_15921_16080# m1_15454_18030# m1_14482_17343# pfet$182
Xpfet$189_5 vdd vdd m1_326_24346# m1_n7513_20152# pfet$189
Xnfet$217_5 m1_26676_16080# m1_26676_16080# vss vss m1_28239_17358# vss nfet$217
Xnfet$195_1 m1_n1263_21786# m1_n1263_21786# m1_354_22513# m1_354_22513# m1_n42_21586#
+ vss nfet$195
Xpfet$187_2 vdd vdd m1_1103_20152# m1_n7401_15478# pfet$187
Xnfet$208_1 m1_28490_22513# m1_28490_22513# vss vss m1_34329_21430# vss nfet$208
Xnfet$222_3 m1_n9336_24346# m1_n9336_24346# vss vss m1_n9854_24542# vss nfet$222
Xpfet$192_0 vdd m1_31535_19792# vdd m1_17939_22513# pfet$192
Xpfet$182_17 vdd vdd m1_n2091_17836# m1_n2250_17343# pfet$182
Xpfet$182_28 vdd m1_2905_18030# vdd m1_1578_16080# pfet$182
Xpfet$182_39 vdd m1_7088_18030# vdd m1_5761_16080# pfet$182
Xpfet$207_3 vdd vdd m1_n4978_24224# vss pfet$207
Xnfet$201_8 m1_n7513_20152# vss m1_26676_16080# vss nfet$201
Xnfet$195_10 m1_19839_21786# m1_19839_21786# m1_21456_22513# m1_21456_22513# m1_21060_21586#
+ vss nfet$195
Xnfet$214_17 m1_21880_15478# m1_21880_15478# m1_n3206_20274# m1_n3206_20274# m1_23924_20470#
+ vss nfet$214
Xnfet$220_0 m1_n3822_20130# m1_n3822_20130# m1_n4485_20152# m1_n4485_20152# m1_n3724_20470#
+ vss nfet$220
Xpfet$205_0 vdd vdd m1_n8625_26174# m1_n9336_24346# pfet$205
Xnfet$199_8 m1_n7383_17599# vss m1_n1133_19550# vss nfet$199
.ends

.subckt asc_drive_buffer$1 vss in vdd out
Xnfet$186_0 out out vss m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# m1_4274_n1060#
+ m1_4274_n1060# out m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# vss vss
+ nfet$186
Xpfet$176_0 vdd vdd m1_3466_n454# in pfet$176
Xpfet$174_0 m1_4274_n1060# vdd vdd m1_4274_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ vdd m1_4002_n1060# m1_4002_n1060# pfet$174
Xnfet$187_0 m1_3466_n454# vss m1_4002_n1060# vss nfet$187
Xnfet$185_0 m1_4274_n1060# vss m1_4002_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ m1_4274_n1060# vss m1_4002_n1060# vss nfet$185
Xpfet$175_0 vdd vdd m1_4002_n1060# m1_3466_n454# pfet$175
Xpfet$173_0 out out m1_4274_n1060# vdd m1_4274_n1060# out vdd vdd m1_4274_n1060# out
+ m1_4274_n1060# m1_4274_n1060# out m1_4274_n1060# vdd m1_4274_n1060# vdd m1_4274_n1060#
+ pfet$173
Xnfet$188_0 in vss m1_3466_n454# vss nfet$188
.ends

.subckt xp_3_1_MUX S0 S1 VDD VSS OUT_1 C_1 B_1 A_1
Xpfet$33_0 VDD A_1 m1_239_n318# m1_n432_458# pfet$33
Xpfet$33_1 VDD C_1 OUT_1 S1 pfet$33
Xpfet$33_2 VDD B_1 m1_239_n318# S0 pfet$33
Xpfet$33_3 VDD m1_239_n318# OUT_1 m1_n432_n1290# pfet$33
Xnfet$39_0 m1_n432_n1290# C_1 OUT_1 VSS nfet$39
Xnfet$39_1 m1_n432_458# B_1 m1_239_n318# VSS nfet$39
Xnfet$39_2 S1 m1_239_n318# OUT_1 VSS nfet$39
Xnfet$39_3 S0 A_1 m1_239_n318# VSS nfet$39
Xpfet$34_0 VDD VDD m1_n432_n1290# S1 pfet$34
Xpfet$34_1 VDD VDD m1_n432_458# S0 pfet$34
Xnfet$40_0 S1 VSS m1_n432_n1290# VSS nfet$40
Xnfet$40_1 S0 VSS m1_n432_458# VSS nfet$40
.ends

.subckt pfet$35 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_954_0# w_n180_n88# a_854_n136#
+ a_n92_0# a_446_n136# a_650_n136# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt nfet$42 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$39 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$45 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt inv1u05u VDD in VSS out
Xpfet$39_0 VDD VDD out in pfet$39
Xnfet$45_0 in VSS out VSS nfet$45
.ends

.subckt pfet$37 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=4.55p ps=15.3u w=7u l=0.5u
.ends

.subckt nfet$43 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$38 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$44 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pass1u05u VDD VSS ind ins clkp clkn
Xpfet$38_0 VDD ind ins clkp pfet$38
Xnfet$44_0 clkn ind ins VSS nfet$44
.ends

.subckt nfet$41 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$40 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.5u
.ends

.subckt nfet$46 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$36 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_954_0# w_n180_n88#
+ a_38_n60# a_n92_0# a_1058_n60# a_854_n60# a_342_0# a_138_0# a_650_n60#
X0 a_954_0# a_854_n60# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n60# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt xp_programmable_basic_pump up vdd s1 s2 s3 s4 down out iref vss
Xpfet$35_18 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$35
Xnfet$42_9 down down vss vss m1_n8807_n11192# vss nfet$42
Xinv1u05u_3 vdd s1 vss inv1u05u_3/out inv1u05u
Xpfet$35_19 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$35
Xnfet$42_10 vss vss vss vss vss vss nfet$42
Xnfet$42_11 vss vss vss vss vss vss nfet$42
Xnfet$42_12 vss vss vss vss vss vss nfet$42
Xnfet$42_13 vss vss vss vss vss vss nfet$42
Xpfet$37_0 vdd vdd vdd vdd pfet$37
Xnfet$43_0 m1_n7879_n12170# pass1u05u_0/ins m1_n7879_n12170# out pass1u05u_0/ins vss
+ nfet$43
Xpfet$37_1 vdd vdd vdd vdd pfet$37
Xpfet$37_2 vdd vdd vdd vdd pfet$37
Xnfet$43_1 m1_n7879_n12170# pass1u05u_0/ins m1_n7879_n12170# out pass1u05u_0/ins vss
+ nfet$43
Xnfet$43_2 vss down vss m1_n7879_n12170# down vss nfet$43
Xpfet$37_3 vdd vdd vdd vdd pfet$37
Xpfet$35_0 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$35
Xpass1u05u_0 vdd vss iref pass1u05u_0/ins inv1u05u_1/out s3 pass1u05u
Xnfet$41_0 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out vss
+ nfet$41
Xnfet$43_3 vss down vss m1_n7879_n12170# down vss nfet$43
Xpfet$35_1 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$35
Xpfet$37_4 vdd vdd vdd vdd pfet$37
Xpass1u05u_1 vdd vss iref pass1u05u_1/ins inv1u05u_2/out s2 pass1u05u
Xnfet$43_4 vss down vss m1_n7879_n12170# down vss nfet$43
Xpfet$37_5 vdd vdd vdd vdd pfet$37
Xpfet$40_0 vdd s3 pass1u05u_5/ins vdd pfet$40
Xnfet$41_1 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out vss
+ nfet$41
Xpfet$35_2 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$35
Xpass1u05u_2 vdd vss iref pass1u05u_2/ins inv1u05u_3/out s1 pass1u05u
Xnfet$41_2 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out vss
+ nfet$41
Xnfet$43_5 vss down vss m1_n7879_n12170# down vss nfet$43
Xpfet$35_3 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$35
Xpfet$37_6 vdd vdd vdd vdd pfet$37
Xpfet$40_1 vdd s2 pass1u05u_4/ins vdd pfet$40
Xnfet$43_6 m1_n7879_n12170# pass1u05u_0/ins m1_n7879_n12170# out pass1u05u_0/ins vss
+ nfet$43
Xpfet$37_7 vdd vdd vdd vdd pfet$37
Xpass1u05u_3 vdd vss pass1u05u_7/ind pass1u05u_3/ins inv1u05u_3/out s1 pass1u05u
Xnfet$41_3 vss vss vss vss vss vss nfet$41
Xpfet$35_4 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$35
Xpfet$40_2 vdd s1 pass1u05u_3/ins vdd pfet$40
Xnfet$43_10 m1_n8607_n8040# pass1u05u_1/ins m1_n8607_n8040# out pass1u05u_1/ins vss
+ nfet$43
Xpass1u05u_4 vdd vss pass1u05u_7/ind pass1u05u_4/ins inv1u05u_2/out s2 pass1u05u
Xnfet$41_4 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out vss
+ nfet$41
Xnfet$43_7 m1_n7879_n12170# pass1u05u_0/ins m1_n7879_n12170# out pass1u05u_0/ins vss
+ nfet$43
Xpfet$35_5 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$35
Xpfet$37_8 vdd vdd vdd vdd pfet$37
Xpfet$40_3 vdd s4 pass1u05u_7/ins vdd pfet$40
Xnfet$43_11 m1_n8144_n9165# iref m1_n8144_n9165# iref iref vss nfet$43
Xnfet$43_8 vss vdd vss m1_n8144_n9165# vdd vss nfet$43
Xpfet$37_9 vdd vdd vdd vdd pfet$37
Xpfet$37_20 vdd vdd vdd vdd pfet$37
Xpass1u05u_5 vdd vss pass1u05u_7/ind pass1u05u_5/ins inv1u05u_1/out s3 pass1u05u
Xnfet$41_5 vss vss vss vss vss vss nfet$41
Xpfet$35_6 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$35
Xnfet$43_12 vss down vss m1_n8607_n8040# down vss nfet$43
Xpfet$37_21 vdd vdd vdd vdd pfet$37
Xpass1u05u_6 vdd vss iref pass1u05u_6/ins inv1u05u_0/out s4 pass1u05u
Xnfet$43_9 m1_n7216_n8262# iref m1_n7216_n8262# pass1u05u_7/ind iref vss nfet$43
Xpfet$37_10 vdd vdd vdd vdd pfet$37
Xnfet$41_6 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out vss
+ nfet$41
Xpfet$35_7 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$35
Xnfet$43_13 vss vdd vss m1_n7216_n8262# vdd vss nfet$43
Xpfet$37_22 vdd vdd vdd vdd pfet$37
Xpass1u05u_7 vdd vss pass1u05u_7/ind pass1u05u_7/ins inv1u05u_0/out s4 pass1u05u
Xnfet$41_7 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out vss
+ nfet$41
Xpfet$35_8 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$35
Xpfet$37_11 vdd vdd vdd vdd pfet$37
Xnfet$43_14 m1_n8607_n8040# pass1u05u_1/ins m1_n8607_n8040# out pass1u05u_1/ins vss
+ nfet$43
Xpfet$37_23 vdd vdd vdd vdd pfet$37
Xnfet$41_8 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out vss
+ nfet$41
Xpfet$35_9 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$35
Xpfet$37_12 vdd vdd vdd vdd pfet$37
Xnfet$43_15 vss down vss m1_n8607_n8040# down vss nfet$43
Xpfet$37_13 vdd vdd vdd vdd pfet$37
Xnfet$41_9 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out vss
+ nfet$41
Xpfet$37_14 vdd vdd vdd vdd pfet$37
Xnfet$46_0 inv1u05u_2/out pass1u05u_1/ins vss vss nfet$46
Xpfet$37_15 vdd vdd vdd vdd pfet$37
Xnfet$46_1 inv1u05u_3/out pass1u05u_2/ins vss vss nfet$46
Xpfet$37_16 vdd vdd vdd vdd pfet$37
Xnfet$46_2 inv1u05u_0/out pass1u05u_6/ins vss vss nfet$46
Xpfet$37_17 vdd vdd vdd vdd pfet$37
Xnfet$46_3 inv1u05u_1/out pass1u05u_0/ins vss vss nfet$46
Xpfet$37_18 vdd vdd vdd vdd pfet$37
Xpfet$37_19 vdd vdd vdd vdd pfet$37
Xnfet$41_10 pass1u05u_2/ins pass1u05u_2/ins m1_n7679_n8960# m1_n7679_n8960# out vss
+ nfet$41
Xpfet$36_0 vdd vdd m1_n4127_3649# vss vss m1_n4127_3649# vdd vss vdd vss vss vdd m1_n4127_3649#
+ vss pfet$36
Xnfet$41_11 vss vss vss vss vss vss nfet$41
Xpfet$35_20 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$35
Xnfet$42_0 down down vss vss m1_n8807_n11192# vss nfet$42
Xpfet$36_1 m1_n5580_883# m1_n5580_883# out pass1u05u_5/ins pass1u05u_5/ins out vdd
+ pass1u05u_5/ins m1_n5580_883# pass1u05u_5/ins pass1u05u_5/ins m1_n5580_883# out
+ pass1u05u_5/ins pfet$36
Xnfet$41_12 down down vss vss m1_n7679_n8960# vss nfet$41
Xnfet$42_1 down down vss vss m1_n8807_n11192# vss nfet$42
Xpfet$36_2 m1_n5580_883# m1_n5580_883# out pass1u05u_5/ins pass1u05u_5/ins out vdd
+ pass1u05u_5/ins m1_n5580_883# pass1u05u_5/ins pass1u05u_5/ins m1_n5580_883# out
+ pass1u05u_5/ins pfet$36
Xpfet$35_21 m1_n6703_2564# m1_n6703_2564# pass1u05u_4/ins out out vdd pass1u05u_4/ins
+ m1_n6703_2564# pass1u05u_4/ins pass1u05u_4/ins m1_n6703_2564# out pass1u05u_4/ins
+ pass1u05u_4/ins pfet$35
Xpfet$35_10 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$35
Xnfet$41_13 vss vss vss vss vss vss nfet$41
Xpfet$35_22 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$35
Xpfet$36_3 m1_n5580_883# m1_n5580_883# out pass1u05u_5/ins pass1u05u_5/ins out vdd
+ pass1u05u_5/ins m1_n5580_883# pass1u05u_5/ins pass1u05u_5/ins m1_n5580_883# out
+ pass1u05u_5/ins pfet$36
Xnfet$42_2 down down vss vss m1_n8807_n11192# vss nfet$42
Xpfet$35_11 vdd vdd up m1_n5450_4559# m1_n5450_4559# vdd up vdd up up vdd m1_n5450_4559#
+ up up pfet$35
Xnfet$41_14 vss vss vss vss vss vss nfet$41
Xpfet$36_4 m1_n5580_883# m1_n5580_883# out pass1u05u_5/ins pass1u05u_5/ins out vdd
+ pass1u05u_5/ins m1_n5580_883# pass1u05u_5/ins pass1u05u_5/ins m1_n5580_883# out
+ pass1u05u_5/ins pfet$36
Xnfet$42_3 down down vss vss m1_n8807_n11192# vss nfet$42
Xpfet$35_23 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$35
Xpfet$35_12 vdd vdd up m1_n6703_2564# m1_n6703_2564# vdd up vdd up up vdd m1_n6703_2564#
+ up up pfet$35
Xnfet$41_15 vss vss vss vss vss vss nfet$41
Xpfet$35_24 m1_n5450_4559# m1_n5450_4559# pass1u05u_3/ins out out vdd pass1u05u_3/ins
+ m1_n5450_4559# pass1u05u_3/ins pass1u05u_3/ins m1_n5450_4559# out pass1u05u_3/ins
+ pass1u05u_3/ins pfet$35
Xpfet$36_5 m1_n4127_3649# m1_n4127_3649# pass1u05u_7/ind pass1u05u_7/ind pass1u05u_7/ind
+ pass1u05u_7/ind vdd pass1u05u_7/ind m1_n4127_3649# pass1u05u_7/ind pass1u05u_7/ind
+ m1_n4127_3649# pass1u05u_7/ind pass1u05u_7/ind pfet$36
Xnfet$42_4 vss vss vss vss vss vss nfet$42
Xpfet$35_13 vdd vdd up m1_n6703_2564# m1_n6703_2564# vdd up vdd up up vdd m1_n6703_2564#
+ up up pfet$35
Xnfet$42_5 vss vss vss vss vss vss nfet$42
Xpfet$35_25 m1_n6703_2564# m1_n6703_2564# pass1u05u_4/ins out out vdd pass1u05u_4/ins
+ m1_n6703_2564# pass1u05u_4/ins pass1u05u_4/ins m1_n6703_2564# out pass1u05u_4/ins
+ pass1u05u_4/ins pfet$35
Xpfet$35_14 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$35
Xnfet$42_6 down down vss vss m1_n8807_n11192# vss nfet$42
Xpfet$35_15 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$35
Xinv1u05u_0 vdd s4 vss inv1u05u_0/out inv1u05u
Xnfet$42_7 down down vss vss m1_n8807_n11192# vss nfet$42
Xpfet$35_16 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$35
Xinv1u05u_1 vdd s3 vss inv1u05u_1/out inv1u05u
Xpfet$35_17 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$35
Xnfet$42_8 down down vss vss m1_n8807_n11192# vss nfet$42
Xinv1u05u_2 vdd s2 vss inv1u05u_2/out inv1u05u
.ends

.subckt asc_hysteresis_buffer$1 vss in vdd out
Xpfet$217_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$217
Xpfet$215_0 vdd vdd m1_884_42# m1_348_648# pfet$215
Xnfet$5_0 m1_1156_42# vss m1_884_42# vss nfet$5
Xnfet$3_0 in vss m1_348_648# vss nfet$3
Xnfet$1_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$1
Xpfet$218_0 vdd vdd m1_884_42# m1_1156_42# pfet$218
Xpfet$216_0 vdd vdd m1_348_648# in pfet$216
Xpfet$214_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd
+ m1_884_42# m1_884_42# pfet$214
Xnfet$4_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$4
Xnfet$2_0 m1_348_648# vss m1_884_42# vss nfet$2
.ends

.subckt pfet$29 a_254_0# a_348_560# w_n180_n88# a_414_0# a_n92_0# a_94_0# a_574_0#
+ a_508_560# a_188_560# a_28_560#
X0 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$35 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt BIAS vdd vss res 200p1 200p2 100n 200n
Xpfet$29_9 vdd res vdd 100n vdd 100n vdd res res res pfet$29
Xpfet$29_10 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$29
Xpfet$29_11 vdd res vdd 200n vdd 200n vdd res res res pfet$29
Xpfet$29_12 vdd res vdd 100n vdd 100n vdd res res res pfet$29
Xpfet$29_13 vdd res vdd res vdd res vdd res res res pfet$29
Xpfet$29_14 vdd res vdd 200n vdd 200n vdd res res res pfet$29
Xpfet$29_15 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$29
Xpfet$29_0 vdd res vdd 200n vdd 200n vdd res res res pfet$29
Xpfet$29_1 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$29
Xnfet$35_0 m1_27_n1423# vss 200p1 m1_27_n1423# vss 200p1 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$35
Xpfet$29_2 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$29
Xnfet$35_1 vss vss vss vss vss vss vss vss vss vss nfet$35
Xpfet$29_3 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$29
Xnfet$35_2 m1_27_n1423# vss 200p2 m1_27_n1423# vss 200p2 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$35
Xpfet$29_5 vdd res vdd 200n vdd 200n vdd res res res pfet$29
Xpfet$29_4 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$29
Xnfet$35_4 m1_27_n1423# vss 200p2 m1_27_n1423# vss 200p2 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$35
Xnfet$35_3 vss vss vss vss vss vss vss vss vss vss nfet$35
Xpfet$29_6 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$29
Xnfet$35_5 m1_27_n1423# vss 200p1 m1_27_n1423# vss 200p1 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$35
Xnfet$35_6 m1_27_n1423# vss m1_27_n1423# m1_27_n1423# vss m1_27_n1423# m1_27_n1423#
+ vss m1_27_n1423# vss nfet$35
Xpfet$29_7 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$29
Xnfet$35_7 m1_27_n1423# vss m1_27_n1423# m1_27_n1423# vss m1_27_n1423# m1_27_n1423#
+ vss m1_27_n1423# vss nfet$35
Xpfet$29_8 vdd res vdd res vdd res vdd res res res pfet$29
.ends

.subckt pfet$18 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$25 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$31 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$23 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$16 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$22 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$21 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt nfet$29 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt pfet$28 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$34 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$27 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$26 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt nfet$32 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt pfet$19 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$25 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$24 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt pfet$17 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$30 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$23 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$22 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$21 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$20 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$28 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$27 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt nfet$33 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt nfet$26 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt nfet$24 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_PFD_DFF_20250831 vss down up vdd fdiv fref
Xpfet$18_2 vdd vdd m1_2068_n5361# m1_2758_n8889# pfet$18
Xpfet$25_3 vdd m1_1452_n8889# m1_2556_n10129# m1_n3884_n9085# pfet$25
Xnfet$31_2 m1_832_n8573# vss m1_1452_n8889# vss nfet$31
Xnfet$31_10 m1_n5867_n10544# vss m1_n5649_n11124# vss nfet$31
Xpfet$23_0 vdd m1_n5428_n3533# vdd m1_n5650_n4045# pfet$23
Xpfet$18_3 vdd vdd m1_1452_n5483# m1_832_n5785# pfet$18
Xpfet$25_4 vdd vdd m1_1452_n8889# m1_832_n8573# pfet$25
Xnfet$31_3 vdd vss m1_1095_n11125# vss nfet$31
Xpfet$16_0 vdd m1_832_n5785# m1_1096_n5165# m1_n3885_n6084# pfet$16
Xpfet$23_1 vdd vdd m1_n5428_n3533# m1_n4678_n3849# pfet$23
Xnfet$31_11 fdiv vss m1_n5867_n10544# vss nfet$31
Xpfet$25_20 vdd m1_n5427_n8573# vdd m1_n5867_n10544# pfet$25
Xpfet$18_4 vdd vdd m1_1095_n4045# vdd pfet$18
Xpfet$25_5 vdd vdd m1_1095_n11125# vdd pfet$25
Xnfet$31_4 m1_n3884_n11124# m1_832_n8573# m1_1096_n9089# vss nfet$31
Xpfet$16_1 vdd m1_1452_n5483# m1_2556_n4049# m1_n3885_n6084# pfet$16
Xnfet$22_0 m1_2068_n5361# m1_2068_n5361# vss vss m1_1550_n5165# vss nfet$22
Xnfet$31_12 m1_n5427_n8573# vss m1_n3884_n9085# vss nfet$31
Xpfet$23_2 vdd m1_n5428_n5842# vdd m1_n5868_n3849# pfet$23
Xpfet$25_10 vdd vdd m1_3349_n9089# m1_2779_n10883# pfet$25
Xpfet$16_2 vdd m1_1095_n4045# m1_832_n5785# m1_n3885_n4045# pfet$16
Xnfet$22_1 m1_1452_n5483# m1_1452_n5483# m1_1096_n5165# m1_1096_n5165# m1_1550_n5165#
+ vss nfet$22
Xpfet$25_6 vdd vdd m1_1096_n9089# m1_1452_n8889# pfet$25
Xnfet$31_5 m1_2758_n8889# vss m1_2068_n8889# vss nfet$31
Xpfet$23_3 vdd vdd m1_n5428_n5842# m1_n4678_n5482# pfet$23
Xpfet$21_0 m1_n1926_n4095# vdd vdd m1_n3099_n4095# pfet$21
Xpfet$25_11 vdd vdd down m1_2779_n10883# pfet$25
Xpfet$25_7 vdd m1_832_n8573# m1_1096_n9089# m1_n3884_n9085# pfet$25
Xnfet$31_6 m1_2779_n10883# vss down vss nfet$31
Xpfet$16_3 vdd m1_2556_n4049# m1_3349_n5165# m1_n3885_n4045# pfet$16
Xnfet$22_2 m1_2556_n4049# m1_2556_n4049# vss vss m1_3015_n4205# vss nfet$22
Xpfet$21_1 m1_n4678_n3849# vdd vdd m1_n1926_n5680# pfet$21
Xpfet$25_12 vdd m1_2556_n10129# m1_3349_n9089# m1_n3884_n11124# pfet$25
Xnfet$22_3 m1_2068_n5361# m1_2068_n5361# m1_2779_n3533# m1_2779_n3533# m1_3015_n4205#
+ vss nfet$22
Xpfet$25_8 vdd m1_1096_n9089# vdd m1_2068_n8889# pfet$25
Xnfet$31_7 m1_2779_n10883# vss m1_3349_n9089# vss nfet$31
Xpfet$21_2 m1_n1926_n5680# vdd vdd m1_n3099_n5680# pfet$21
Xpfet$25_13 vdd vdd m1_n5427_n8573# m1_n4677_n8889# pfet$25
Xpfet$25_9 vdd vdd m1_2068_n8889# m1_2758_n8889# pfet$25
Xnfet$31_8 m1_n3884_n9085# m1_2556_n10129# m1_3349_n9089# vss nfet$31
Xpfet$21_3 m1_n4678_n5482# vdd vdd m1_n1926_n4095# pfet$21
Xpfet$25_14 vdd vdd m1_n3884_n11124# m1_n5427_n10882# pfet$25
Xnfet$31_9 m1_n5427_n10882# vss m1_n3884_n11124# vss nfet$31
Xpfet$25_15 vdd m1_n5427_n10882# vdd m1_n5649_n11124# pfet$25
Xpfet$25_16 vdd vdd m1_n5427_n10882# m1_n4677_n10522# pfet$25
Xnfet$29_0 m1_n3885_n4045# vss m1_n3099_n4095# vss nfet$29
Xpfet$25_17 vdd vdd m1_n5649_n11124# m1_n5867_n10544# pfet$25
Xpfet$28_0 vdd m1_5895_n8089# vdd down pfet$28
Xnfet$29_1 m1_n3885_n6084# vss m1_n3099_n5680# vss nfet$29
Xpfet$25_18 vdd vdd m1_n5867_n10544# fdiv pfet$25
Xnfet$34_0 up up m1_5895_n8089# m1_5895_n8089# m1_5043_n9245# vss nfet$34
Xpfet$28_1 vdd vdd m1_5895_n8089# up pfet$28
Xpfet$25_19 vdd vdd m1_n3884_n9085# m1_n5427_n8573# pfet$25
Xnfet$34_1 down down vss vss m1_5043_n9245# vss nfet$34
Xnfet$27_0 m1_n5428_n3533# vss m1_n3885_n4045# vss nfet$27
Xnfet$27_1 m1_n5868_n3849# vss m1_n5650_n4045# vss nfet$27
Xpfet$26_0 vdd vdd m1_n3098_n10720# m1_n3884_n11124# pfet$26
Xnfet$32_0 m1_n3884_n11124# vss m1_n3098_n10720# vss nfet$32
Xpfet$26_1 vdd vdd m1_n3098_n9135# m1_n3884_n9085# pfet$26
Xnfet$27_2 m1_n5428_n5842# vss m1_n3885_n6084# vss nfet$27
Xpfet$19_0 vdd vdd m1_2758_n8889# m1_4978_n5483# pfet$19
Xnfet$27_3 fref vss m1_n5868_n3849# vss nfet$27
Xnfet$32_1 m1_n3884_n9085# vss m1_n3098_n9135# vss nfet$32
Xnfet$25_0 m1_5895_n8089# vss m1_5464_n5483# vss nfet$25
Xnfet$25_1 m1_5464_n5483# vss m1_4978_n5483# vss nfet$25
Xpfet$24_0 vdd vdd m1_n3099_n4095# m1_n3885_n4045# pfet$24
Xpfet$17_0 vdd vdd m1_1096_n5165# m1_1452_n5483# pfet$17
Xnfet$30_0 m1_2556_n10129# m1_2556_n10129# vss vss m1_3015_n10205# vss nfet$30
Xpfet$24_1 vdd vdd m1_n3099_n5680# m1_n3885_n6084# pfet$24
Xpfet$17_1 vdd m1_1096_n5165# vdd m1_2068_n5361# pfet$17
Xnfet$30_1 m1_1452_n8889# m1_1452_n8889# m1_1096_n9089# m1_1096_n9089# m1_1550_n9245#
+ vss nfet$30
Xnfet$23_0 m1_2779_n3533# vss up vss nfet$23
Xpfet$17_2 vdd m1_2779_n3533# vdd m1_2556_n4049# pfet$17
Xnfet$30_2 m1_2068_n8889# m1_2068_n8889# vss vss m1_1550_n9245# vss nfet$30
Xpfet$22_0 vdd vdd m1_n3885_n4045# m1_n5428_n3533# pfet$22
Xnfet$23_1 m1_2779_n3533# vss m1_3349_n5165# vss nfet$23
Xpfet$17_3 vdd vdd m1_2779_n3533# m1_2068_n5361# pfet$17
Xnfet$23_2 m1_2758_n8889# vss m1_2068_n5361# vss nfet$23
Xnfet$30_3 m1_2068_n8889# m1_2068_n8889# m1_2779_n10883# m1_2779_n10883# m1_3015_n10205#
+ vss nfet$30
Xpfet$22_1 vdd vdd m1_n5650_n4045# m1_n5868_n3849# pfet$22
Xnfet$23_3 m1_832_n5785# vss m1_1452_n5483# vss nfet$23
Xnfet$21_0 m1_n3885_n4045# m1_832_n5785# m1_1096_n5165# vss nfet$21
Xnfet$30_4 m1_n4677_n10522# m1_n4677_n10522# m1_n5427_n10882# m1_n5427_n10882# m1_n5191_n10204#
+ vss nfet$30
Xpfet$22_2 vdd vdd m1_n3885_n6084# m1_n5428_n5842# pfet$22
Xnfet$23_4 vdd vss m1_1095_n4045# vss nfet$23
Xnfet$30_5 m1_n5649_n11124# m1_n5649_n11124# vss vss m1_n5191_n10204# vss nfet$30
Xnfet$21_1 m1_n3885_n4045# m1_1452_n5483# m1_2556_n4049# vss nfet$21
Xpfet$22_3 vdd vdd m1_n5868_n3849# fref pfet$22
Xpfet$20_0 vdd vdd m1_5464_n5483# m1_5895_n8089# pfet$20
Xnfet$21_2 m1_n3885_n6084# m1_1095_n4045# m1_832_n5785# vss nfet$21
Xnfet$30_6 m1_n4677_n8889# m1_n4677_n8889# m1_n5427_n8573# m1_n5427_n8573# m1_n5191_n9245#
+ vss nfet$30
Xpfet$20_1 vdd vdd m1_4978_n5483# m1_5464_n5483# pfet$20
Xnfet$30_7 m1_n5867_n10544# m1_n5867_n10544# vss vss m1_n5191_n9245# vss nfet$30
Xnfet$21_3 m1_n3885_n6084# m1_2556_n4049# m1_3349_n5165# vss nfet$21
Xnfet$28_0 m1_n4678_n3849# m1_n4678_n3849# m1_n5428_n3533# m1_n5428_n3533# m1_n5192_n4205#
+ vss nfet$28
Xnfet$28_1 m1_n5650_n4045# m1_n5650_n4045# vss vss m1_n5192_n4205# vss nfet$28
Xpfet$27_0 m1_n4677_n8889# vdd vdd m1_n1925_n10720# pfet$27
Xpfet$27_1 m1_n1925_n10720# vdd vdd m1_n3098_n10720# pfet$27
Xnfet$28_2 m1_n4678_n5482# m1_n4678_n5482# m1_n5428_n5842# m1_n5428_n5842# m1_n5192_n5164#
+ vss nfet$28
Xnfet$33_0 m1_n4677_n8889# m1_n1925_n10720# vss vss nfet$33
Xnfet$28_3 m1_n5868_n3849# m1_n5868_n3849# vss vss m1_n5192_n5164# vss nfet$28
Xnfet$33_1 m1_n1925_n10720# m1_n3098_n10720# vss vss nfet$33
Xpfet$27_2 m1_n4677_n10522# vdd vdd m1_n1925_n9135# pfet$27
Xnfet$26_0 m1_n1926_n4095# m1_n3099_n4095# vss vss nfet$26
Xpfet$25_0 vdd vdd m1_2779_n10883# m1_2068_n8889# pfet$25
Xnfet$33_2 m1_n4677_n10522# m1_n1925_n9135# vss vss nfet$33
Xpfet$27_3 m1_n1925_n9135# vdd vdd m1_n3098_n9135# pfet$27
Xnfet$26_1 m1_n4678_n3849# m1_n1926_n5680# vss vss nfet$26
Xnfet$33_3 m1_n1925_n9135# m1_n3098_n9135# vss vss nfet$33
Xnfet$26_2 m1_n1926_n5680# m1_n3099_n5680# vss vss nfet$26
Xpfet$25_1 vdd m1_2779_n10883# vdd m1_2556_n10129# pfet$25
Xnfet$31_0 m1_n3884_n9085# m1_1095_n11125# m1_832_n8573# vss nfet$31
Xpfet$18_0 vdd vdd m1_3349_n5165# m1_2779_n3533# pfet$18
Xpfet$25_2 vdd m1_1095_n11125# m1_832_n8573# m1_n3884_n11124# pfet$25
Xnfet$31_1 m1_n3884_n11124# m1_1452_n8889# m1_2556_n10129# vss nfet$31
Xnfet$26_3 m1_n4678_n5482# m1_n1926_n4095# vss vss nfet$26
Xnfet$24_0 m1_4978_n5483# vss m1_2758_n8889# vss nfet$24
Xpfet$18_1 vdd vdd up m1_2779_n3533# pfet$18
.ends

.subckt pfet$30 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=9.75p pd=31.3u as=9.75p ps=31.3u w=15u l=0.5u
.ends

.subckt nfet$38 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$36 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.5u
.ends

.subckt cap_mim m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
.ends

.subckt pfet$31 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=9.75p pd=31.3u as=9.75p ps=31.3u w=15u l=0.5u
.ends

.subckt nfet$37 a_n84_0# a_38_n132# a_138_0# VSUBS
X0 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.5u
.ends

.subckt pfet$32 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt CSRVCO_20250823 vctrl vosc vdd vss
Xpfet$30_0 vdd vdd m1_n12264_2422# m1_n16019_266# pfet$30
Xpfet$30_1 vdd vdd m1_n14208_3657# m1_n16019_266# pfet$30
Xpfet$30_2 vdd vdd m1_n13722_3340# m1_n16019_266# pfet$30
Xpfet$30_3 vdd m1_n16019_266# vdd m1_n16019_266# pfet$30
Xpfet$30_10 vdd m1_n14208_3657# m1_n10810_266# m1_n11296_266# pfet$30
Xpfet$30_4 vdd vdd m1_n13236_3035# m1_n16019_266# pfet$30
Xpfet$30_11 vdd m1_n12264_2422# m1_n11916_1270# m1_n9352_266# pfet$30
Xpfet$30_12 vdd m1_n14693_3963# m1_n11296_266# m1_n11782_266# pfet$30
Xpfet$30_5 vdd vdd m1_n14693_3963# m1_n16019_266# pfet$30
Xpfet$30_13 vdd m1_n13722_3340# m1_n10324_266# m1_n10810_266# pfet$30
Xpfet$30_6 vdd vdd m1_n12750_2729# m1_n16019_266# pfet$30
Xnfet$38_0 m1_n8380_274# vss vosc vss nfet$38
Xpfet$30_14 vdd m1_n15180_4275# m1_n11782_266# m1_n11916_1270# pfet$30
Xpfet$30_7 vdd vdd m1_n15180_4275# m1_n16019_266# pfet$30
Xnfet$38_1 m1_n11916_1270# vss m1_n8380_274# vss nfet$38
Xpfet$30_8 vdd m1_n13236_3035# m1_n9838_266# m1_n10324_266# pfet$30
Xpfet$30_9 vdd m1_n12750_2729# m1_n9352_266# m1_n9838_266# pfet$30
Xnfet$36_0 m1_n9838_266# m1_n12754_674# m1_n9352_266# vss nfet$36
Xcap_mim_0 vss m1_n11296_266# cap_mim
Xnfet$36_1 vctrl vss m1_n12268_985# vss nfet$36
Xcap_mim_1 vss m1_n10810_266# cap_mim
Xnfet$36_2 vctrl vss m1_n14283_186# vss nfet$36
Xcap_mim_2 vss m1_n10324_266# cap_mim
Xnfet$36_3 vctrl vss m1_n13794_186# vss nfet$36
Xnfet$36_4 vctrl vss m1_n13240_368# vss nfet$36
Xcap_mim_3 vss m1_n11916_1270# cap_mim
Xcap_mim_5 vss m1_n9838_266# cap_mim
Xnfet$36_5 vctrl vss m1_n12754_674# vss nfet$36
Xcap_mim_4 vss m1_n9352_266# cap_mim
Xcap_mim_6 vss m1_n11782_266# cap_mim
Xnfet$36_6 vctrl m1_n16019_266# vss vss nfet$36
Xpfet$31_0 vdd vdd vdd vdd pfet$31
Xnfet$36_7 vctrl vss m1_n15245_186# vss nfet$36
Xpfet$31_1 vdd vdd vdd vdd pfet$31
Xnfet$36_9 m1_n10324_266# m1_n13240_368# m1_n9838_266# vss nfet$36
Xnfet$36_8 vctrl vss m1_n14765_186# vss nfet$36
Xnfet$37_0 vss vss vss vss nfet$37
Xnfet$37_1 vss vss vss vss nfet$37
Xnfet$36_10 m1_n9352_266# m1_n12268_985# m1_n11916_1270# vss nfet$36
Xnfet$36_11 m1_n11916_1270# m1_n15245_186# m1_n11782_266# vss nfet$36
Xnfet$36_12 m1_n11782_266# m1_n14765_186# m1_n11296_266# vss nfet$36
Xnfet$36_13 m1_n11296_266# m1_n14283_186# m1_n10810_266# vss nfet$36
Xnfet$36_14 m1_n10810_266# m1_n13794_186# m1_n10324_266# vss nfet$36
Xpfet$32_0 vdd vdd vosc m1_n8380_274# pfet$32
Xpfet$32_1 vdd vdd m1_n8380_274# m1_n11916_1270# pfet$32
.ends

.subckt top_level_20250912_nosc vdd vss i_cp_100u div_def div_prc_s8 div_prc_s7 div_prc_s6
+ div_prc_s5 div_prc_s4 div_prc_s3 div_prc_s2 div_prc_s1 div_prc_s0 div_out div_in
+ div_swc_s0 div_swc_s1 div_swc_s2 div_swc_s3 div_swc_s4 div_swc_s5 div_swc_s6 div_swc_s7
+ div_swc_s8 lock ref ext_pfd_div ext_pfd_ref ext_pfd_up ext_pfd_down mx_pfd_s1 mx_pfd_s0
+ up down cp_s1 cp_s2 cp_s3 cp_s4 filter_in out filter_out ext_vco_in ext_vco_out
+ mx_vco_s0 mx_vco_s1 div_rpc_s0 div_rsc_s0 div_rsc_s1 div_rpc_s1 div_rsc_s2 div_rpc_s2
+ div_rsc_s3 div_rsc_s4 div_rsc_s5 div_rsc_s6 div_rsc_s7 div_rsc_s8 div_rpc_s3 div_rpc_s4
+ div_rpc_s5 div_rpc_s6 div_rpc_s7 div_rpc_s8 mx_ref_s1 mx_ref_s0
Xasc_drive_buffer_up_0 vss asc_drive_buffer_up_0/out xp_3_1_MUX_2/OUT_1 vdd asc_drive_buffer_up
Xasc_dual_psd_def_20250809_0 vdd vss div_prc_s0 div_prc_s1 div_prc_s2 div_prc_s3 div_prc_s4
+ div_prc_s5 div_prc_s6 div_prc_s7 div_prc_s8 xp_3_1_MUX_4/OUT_1 div_swc_s0 div_swc_s1
+ div_swc_s2 div_swc_s3 div_swc_s4 div_swc_s5 div_swc_s6 div_swc_s7 div_swc_s8 asc_drive_buffer_0/in
+ div_def asc_dual_psd_def_20250809
Xasc_drive_buffer_0 vss asc_drive_buffer_0/in vdd div_in asc_drive_buffer
Xxp_3_1_MUX$1_0 mx_ref_s0 mx_ref_s1 vdd vss xp_3_1_MUX$1_0/OUT_1 xp_3_1_MUX$1_1/C_1
+ xp_3_1_MUX$1_0/B_1 xp_3_1_MUX$1_0/A_1 xp_3_1_MUX$1
Xasc_drive_buffer_1 vss xp_3_1_MUX_0/OUT_1 vdd out asc_drive_buffer
Xxp_3_1_MUX$1_1 mx_ref_s0 mx_ref_s1 vdd vss xp_3_1_MUX$1_1/OUT_1 xp_3_1_MUX$1_1/C_1
+ xp_3_1_MUX$1_1/B_1 xp_3_1_MUX$1_1/A_1 xp_3_1_MUX$1
Xasc_drive_buffer_2 vss xp_3_1_MUX_4/OUT_1 vdd div_out asc_drive_buffer
Xasc_drive_buffer_3 vss asc_drive_buffer_3/in vdd lock asc_drive_buffer
Xasc_hysteresis_buffer_0 vss xp_3_1_MUX$1_1/OUT_1 vdd xp_3_1_MUX_3/OUT_1 asc_hysteresis_buffer
Xasc_drive_buffer_4 vss xp_3_1_MUX_2/OUT_1 vdd up asc_drive_buffer
Xasc_lock_detector_20250826_0 xp_3_1_MUX_3/OUT_1 vdd xp_3_1_MUX_4/OUT_1 asc_drive_buffer_3/in
+ vss asc_lock_detector_20250826
Xasc_drive_buffer_5 vss xp_3_1_MUX_5/OUT_1 vdd down asc_drive_buffer
Xasc_drive_buffer_6 vss xp_3_1_MUX_5/OUT_1 vdd asc_drive_buffer_6/out asc_drive_buffer
Xasc_dual_psd_def_20250809$1_0 vdd vss div_rpc_s0 div_rpc_s1 div_rpc_s2 div_rpc_s3
+ div_rpc_s4 div_rpc_s5 div_rpc_s6 div_rpc_s7 div_rpc_s8 xp_3_1_MUX$1_1/B_1 div_rsc_s0
+ div_rsc_s1 div_rsc_s2 div_rsc_s3 div_rsc_s4 div_rsc_s5 div_rsc_s6 div_rsc_s7 div_rsc_s8
+ xp_3_1_MUX$1_0/B_1 vss asc_dual_psd_def_20250809$1
Xasc_drive_buffer$1_0 vss xp_3_1_MUX_0/OUT_1 vdd asc_drive_buffer_0/in asc_drive_buffer$1
Xxp_3_1_MUX_0 mx_vco_s0 mx_vco_s1 vdd vss xp_3_1_MUX_0/OUT_1 xp_3_1_MUX_0/C_1 xp_3_1_MUX_0/B_1
+ ext_vco_out xp_3_1_MUX
Xxp_3_1_MUX_1 mx_vco_s0 mx_vco_s1 vdd vss filter_out xp_3_1_MUX_1/C_1 xp_3_1_MUX_1/B_1
+ ext_vco_in xp_3_1_MUX
Xxp_3_1_MUX_2 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX_2/OUT_1 xp_3_1_MUX_2/C_1 xp_3_1_MUX_2/B_1
+ ext_pfd_up xp_3_1_MUX
Xxp_3_1_MUX_3 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX_3/OUT_1 xp_3_1_MUX_3/C_1 xp_3_1_MUX_3/B_1
+ ext_pfd_ref xp_3_1_MUX
Xxp_3_1_MUX_4 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX_4/OUT_1 xp_3_1_MUX_4/C_1 xp_3_1_MUX_4/B_1
+ ext_pfd_div xp_3_1_MUX
Xxp_3_1_MUX_5 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX_5/OUT_1 xp_3_1_MUX_5/C_1 xp_3_1_MUX_5/B_1
+ ext_pfd_down xp_3_1_MUX
Xxp_programmable_basic_pump_0 asc_drive_buffer_up_0/out vdd cp_s1 cp_s2 cp_s3 cp_s4
+ asc_drive_buffer_6/out filter_in BIAS_0/100n vss xp_programmable_basic_pump
Xasc_hysteresis_buffer$1_0 vss ref vdd xp_3_1_MUX$1_0/OUT_1 asc_hysteresis_buffer$1
XBIAS_0 vdd vss i_cp_100u BIAS_0/200p1 BIAS_0/200p2 BIAS_0/100n BIAS_0/200n BIAS
Xasc_PFD_DFF_20250831_0 vss xp_3_1_MUX_5/C_1 xp_3_1_MUX_2/C_1 vdd xp_3_1_MUX_4/C_1
+ xp_3_1_MUX_3/C_1 asc_PFD_DFF_20250831
Xasc_PFD_DFF_20250831_1 vss xp_3_1_MUX_2/B_1 xp_3_1_MUX_5/B_1 vdd xp_3_1_MUX_4/B_1
+ xp_3_1_MUX_3/B_1 asc_PFD_DFF_20250831
XCSRVCO_20250823_0 xp_3_1_MUX_1/C_1 xp_3_1_MUX_0/C_1 vdd vss CSRVCO_20250823
.ends

