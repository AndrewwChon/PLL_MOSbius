* Extracted by KLayout with GF180MCU LVS runset on : 29/07/2025 06:12

.SUBCKT asc_NAND VSS B A VDD
M$1 VDD B \$4 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$2 \$4 A VDD VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$3 \$3 B VSS VSS nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$4 \$4 A \$3 VSS nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
.ENDS asc_NAND
