* Extracted by KLayout with GF180MCU LVS runset on : 08/08/2025 02:56

.SUBCKT asc_XNOR VSS VDD A B OUT
M$1 VDD A \$7 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$2 VDD B \$9 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$3 \$19 \$9 OUT VDD pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U PD=13.3U
M$4 \$26 A VDD VDD pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U PD=13.3U
M$5 OUT B \$26 VDD pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U PD=13.3U
M$6 VDD \$7 \$19 VDD pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U PD=13.3U
M$7 VSS A \$7 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$8 \$5 \$9 VSS VSS nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$9 OUT A \$5 VSS nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$10 \$6 B VSS VSS nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$11 OUT \$7 \$6 VSS nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$12 VSS B \$9 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
.ENDS asc_XNOR
