** sch_path: /foss/designs/switch_matrix_gf180mcu_9t5v0-main/DFF_flatten/DFF_flatten.sch
.subckt DFF_flatten D Q PHI_1 PHI_2 VDDd VSSd
*.PININFO D:I PHI_1:I PHI_2:I Q:O VDDd:B VSSd:B
* noconn VSSd
* noconn VDDd
xmain D PHI_1 out_m VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1
xsecondary out_m PHI_2 Q VDDd VDDd VSSd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1
.ends
