* Extracted by KLayout with GF180MCU LVS runset on : 05/09/2025 03:59

.SUBCKT qw_NOLclk PHI_1 VSSd PHI_2 CLK VDDd
M$1 \$2 \$11 VDDd VDDd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$2 VDDd \$2 \$3 VDDd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$3 \$3 \$1 VDDd VDDd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$4 PHI_1 \$3 VDDd VDDd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$5 \$12 PHI_1 VDDd VDDd pfet_03v3 L=2U W=1U AS=0.65P AD=0.65P PS=3.3U PD=3.3U
M$6 \$13 \$12 VDDd VDDd pfet_03v3 L=4U W=1U AS=0.65P AD=0.65P PS=3.3U PD=3.3U
M$7 \$52 \$13 VDDd VDDd pfet_03v3 L=4U W=1U AS=0.65P AD=0.65P PS=3.3U PD=3.3U
M$8 \$46 PHI_2 VDDd VDDd pfet_03v3 L=2U W=1U AS=0.65P AD=0.65P PS=3.3U PD=3.3U
M$9 \$47 \$46 VDDd VDDd pfet_03v3 L=4U W=1U AS=0.65P AD=0.65P PS=3.3U PD=3.3U
M$10 \$1 \$47 VDDd VDDd pfet_03v3 L=4U W=1U AS=0.65P AD=0.65P PS=3.3U PD=3.3U
M$11 \$11 CLK VDDd VDDd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$12 VDDd \$11 \$44 VDDd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$13 \$44 \$52 VDDd VDDd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$14 PHI_2 \$44 VDDd VDDd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$15 \$2 \$11 VSSd VSSd nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$16 \$23 \$2 VSSd VSSd nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$18 \$23 \$1 \$3 VSSd nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U PD=4.74U
M$20 PHI_1 \$3 VSSd VSSd nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$21 \$12 PHI_1 VSSd VSSd nfet_03v3 L=2U W=0.5U AS=0.305P AD=0.305P PS=2.22U
+ PD=2.22U
M$22 \$13 \$12 VSSd VSSd nfet_03v3 L=4U W=0.5U AS=0.305P AD=0.305P PS=2.22U
+ PD=2.22U
M$23 \$52 \$13 VSSd VSSd nfet_03v3 L=4U W=0.5U AS=0.305P AD=0.305P PS=2.22U
+ PD=2.22U
M$24 \$46 PHI_2 VSSd VSSd nfet_03v3 L=2U W=0.5U AS=0.305P AD=0.305P PS=2.22U
+ PD=2.22U
M$25 \$47 \$46 VSSd VSSd nfet_03v3 L=4U W=0.5U AS=0.305P AD=0.305P PS=2.22U
+ PD=2.22U
M$26 \$1 \$47 VSSd VSSd nfet_03v3 L=4U W=0.5U AS=0.305P AD=0.305P PS=2.22U
+ PD=2.22U
M$27 \$11 CLK VSSd VSSd nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$28 \$31 \$11 VSSd VSSd nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$30 \$31 \$52 \$44 VSSd nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$32 PHI_2 \$44 VSSd VSSd nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
.ENDS qw_NOLclk
