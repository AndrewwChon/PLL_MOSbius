* Extracted by KLayout with GF180MCU LVS runset on : 09/09/2025 21:45

.SUBCKT asc_dual_psd_def_20250809 vdd sd9 sd8 sd7 sd6 sd5 sd4 sd3 sd2 sd1 vss
+ fout define fin pd1 pd2 pd3 pd4 pd5 pd6 pd7 pd8 pd9
M$1 vdd sd9 \$77 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$2 vdd \$119 \$78 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$3 \$78 \$120 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$4 \$79 \$3 \$120 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$5 vdd \$121 \$79 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$6 \$81 \$80 \$121 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$7 vdd \$78 \$81 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$8 vdd \$3 \$80 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$9 vdd sd8 \$4 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$10 vdd \$123 \$82 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$11 \$82 \$124 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$12 \$83 \$5 \$124 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$13 vdd \$125 \$83 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$14 \$85 \$84 \$125 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$15 vdd \$82 \$85 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$16 vdd \$5 \$84 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$17 vdd sd7 \$86 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$18 vdd \$127 \$87 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$19 \$87 \$128 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$20 \$88 \$6 \$128 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$21 vdd \$129 \$88 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$22 \$90 \$89 \$129 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$23 vdd \$87 \$90 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$24 vdd \$6 \$89 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$25 vdd sd6 \$91 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$26 vdd \$454 \$131 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$27 \$131 \$132 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$28 \$92 \$7 \$132 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$29 vdd \$133 \$92 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$30 \$94 \$93 \$133 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$31 vdd \$131 \$94 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$32 vdd \$7 \$93 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$33 vdd sd5 \$8 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$34 vdd \$458 \$135 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$35 \$135 \$136 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$36 \$95 \$9 \$136 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$37 vdd \$137 \$95 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$38 \$97 \$96 \$137 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$39 vdd \$135 \$97 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$40 vdd \$9 \$96 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$41 vdd sd4 \$98 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$42 vdd \$139 \$99 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$43 \$99 \$140 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$44 \$100 \$10 \$140 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$45 vdd \$141 \$100 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$46 \$102 \$101 \$141 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$47 vdd \$99 \$102 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$48 vdd \$10 \$101 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$49 vdd sd3 \$103 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$50 vdd \$143 \$104 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$51 \$104 \$144 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$52 \$105 \$11 \$144 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$53 vdd \$145 \$105 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$54 \$107 \$106 \$145 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$55 vdd \$104 \$107 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$56 vdd \$11 \$106 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$57 vdd sd2 \$108 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$58 vdd \$468 \$109 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$59 \$109 \$147 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$60 \$110 \$12 \$147 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$61 vdd \$148 \$110 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$62 \$112 \$111 \$148 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$63 vdd \$109 \$112 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$64 vdd \$12 \$111 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$65 vdd sd1 \$113 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$66 vdd \$150 \$114 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$67 \$114 \$151 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$68 \$115 \$13 \$151 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$69 vdd \$152 \$115 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$70 \$117 \$116 \$152 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$71 vdd \$114 \$117 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$72 vdd \$13 \$116 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$73 vdd \$78 \$443 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$74 \$444 \$78 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$75 \$120 \$80 \$444 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$76 \$119 \$1 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$77 vdd \$119 \$445 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$78 \$445 \$79 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$79 \$121 \$3 \$445 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$80 vdd \$446 \$3 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$81 vdd \$82 \$446 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$82 \$447 \$82 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$83 \$124 \$84 \$447 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$84 \$123 \$1 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$85 vdd \$123 \$448 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$86 \$448 \$83 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$87 \$125 \$5 \$448 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$88 vdd \$449 \$5 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$89 vdd \$87 \$449 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$90 \$450 \$87 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$91 \$128 \$89 \$450 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$92 \$127 \$1 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$93 vdd \$127 \$451 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$94 \$451 \$88 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$95 \$129 \$6 \$451 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$96 vdd \$452 \$6 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$97 vdd \$131 \$452 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$98 \$453 \$131 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$99 \$132 \$93 \$453 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$100 \$454 \$1 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$101 vdd \$454 \$455 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$102 \$455 \$92 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$103 \$133 \$7 \$455 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$104 vdd \$456 \$7 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$105 vdd \$135 \$456 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$106 \$457 \$135 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$107 \$136 \$96 \$457 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$108 \$458 \$1 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$109 vdd \$458 \$459 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$110 \$459 \$95 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$111 \$137 \$9 \$459 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$112 vdd \$460 \$9 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$113 vdd \$99 \$460 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$114 \$461 \$99 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$115 \$140 \$101 \$461 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$116 \$139 \$1 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$117 vdd \$139 \$462 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$118 \$462 \$100 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$119 \$141 \$10 \$462 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$120 vdd \$463 \$10 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$121 vdd \$104 \$463 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$122 \$464 \$104 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$123 \$144 \$106 \$464 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$124 \$143 \$1 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$125 vdd \$143 \$465 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$126 \$465 \$105 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$127 \$145 \$11 \$465 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$128 vdd \$466 \$11 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$129 vdd \$109 \$466 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$130 \$467 \$109 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$131 \$147 \$111 \$467 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$132 \$468 \$1 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$133 vdd \$468 \$469 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$134 \$469 \$110 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$135 \$148 \$12 \$469 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$136 vdd \$470 \$12 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$137 vdd \$114 \$470 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$138 \$471 \$114 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$139 \$151 \$116 \$471 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$140 \$150 \$1 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$141 vdd \$150 \$472 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$142 \$472 \$115 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$143 \$152 \$13 \$472 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$144 vdd \$473 \$13 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$145 \$739 \$788 \$738 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$147 \$739 \$1 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$149 vdd \$741 \$740 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$150 vdd \$789 \$741 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$151 \$741 \$681 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$152 \$743 \$745 \$742 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$154 \$743 \$744 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$156 vdd \$689 \$744 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$157 \$744 \$688 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$158 vdd \$687 \$745 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$159 \$745 \$686 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$160 \$746 \$443 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$161 \$747 \$746 \$681 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$163 \$748 \$443 \$681 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$165 \$748 \$77 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$167 \$747 \$749 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$169 vdd \$77 \$749 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$170 \$750 \$446 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$171 \$751 \$750 \$682 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$173 \$752 \$446 \$682 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$175 \$752 \$4 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$177 \$751 \$753 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$179 vdd \$4 \$753 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$180 \$754 \$449 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$181 \$755 \$754 \$683 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$183 \$756 \$449 \$683 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$185 \$756 \$86 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$187 \$755 \$757 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$189 vdd \$86 \$757 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$190 \$758 \$452 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$191 \$759 \$758 \$684 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$193 \$760 \$452 \$684 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$195 \$760 \$91 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$197 \$759 \$761 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$199 vdd \$91 \$761 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$200 \$762 \$456 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$201 \$763 \$762 \$685 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$203 \$764 \$456 \$685 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$205 \$764 \$8 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$207 \$763 \$765 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$209 vdd \$8 \$765 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$210 \$766 \$460 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$211 \$767 \$766 \$686 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$213 \$768 \$460 \$686 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$215 \$768 \$98 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$217 \$767 \$769 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$219 vdd \$98 \$769 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$220 \$770 \$463 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$221 \$771 \$770 \$687 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$223 \$772 \$463 \$687 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$225 \$772 \$103 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$227 \$771 \$773 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$229 vdd \$103 \$773 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$230 \$774 \$466 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$231 \$775 \$774 \$688 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$233 \$776 \$466 \$688 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$235 \$776 \$108 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$237 \$775 \$777 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$239 vdd \$108 \$777 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$240 \$778 \$470 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$241 \$779 \$778 \$689 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$243 \$780 \$470 \$689 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$245 \$780 \$113 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$247 \$779 \$781 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$249 vdd \$113 \$781 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$250 vdd \$1033 \$782 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$251 \$782 \$1031 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$252 vdd \$1029 \$783 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$253 \$783 \$1027 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$254 \$784 \$783 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$256 \$784 \$782 \$785 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$258 vdd \$785 \$786 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$259 \$786 \$866 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$260 \$787 \$786 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$261 vdd \$790 \$1 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$262 \$1217 \$740 \$788 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$264 \$1217 \$738 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$266 vdd \$1088 \$789 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$267 vdd \$742 \$1088 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$268 \$1088 \$1089 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$269 \$1218 \$1016 \$1089 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$271 \$1218 \$1090 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$273 vdd \$685 \$1090 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$274 \$1090 \$684 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$275 vdd \$683 \$1016 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$276 \$1016 \$682 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$277 \$1092 \$1091 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$278 \$1219 \$1092 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$280 \$1220 \$1091 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$282 \$1220 \$1094 \$1019 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$284 \$1219 \$1095 \$1019 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$286 vdd \$1094 \$1095 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$287 \$1097 \$1096 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$288 \$1221 \$1097 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$290 \$1222 \$1096 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$292 \$1222 \$1099 \$1021 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$294 \$1221 \$1100 \$1021 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$296 vdd \$1099 \$1100 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$297 \$1102 \$1101 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$298 \$1223 \$1102 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$300 \$1224 \$1101 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$302 \$1224 \$1104 \$1023 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$304 \$1223 \$1105 \$1023 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$306 vdd \$1104 \$1105 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$307 \$1107 \$1106 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$308 \$1225 \$1107 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$310 \$1226 \$1106 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$312 \$1226 \$1109 \$1025 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$314 \$1225 \$1110 \$1025 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$316 vdd \$1109 \$1110 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$317 \$1112 \$1111 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$318 \$1227 \$1112 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$320 \$1228 \$1111 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$322 \$1228 \$1114 \$1027 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$324 \$1227 \$1115 \$1027 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$326 vdd \$1114 \$1115 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$327 \$1117 \$1116 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$328 \$1229 \$1117 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$330 \$1230 \$1116 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$332 \$1230 \$1119 \$1029 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$334 \$1229 \$1120 \$1029 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$336 vdd \$1119 \$1120 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$337 \$1122 \$1121 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$338 \$1231 \$1122 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$340 \$1232 \$1121 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$342 \$1232 \$1124 \$1031 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$344 \$1231 \$1125 \$1031 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$346 vdd \$1124 \$1125 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$347 \$1127 \$1126 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$348 \$1233 \$1127 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$350 \$1234 \$1126 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$352 \$1234 \$1129 \$1033 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$354 \$1233 \$1130 \$1033 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$356 vdd \$1129 \$1130 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$357 \$1132 \$1131 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$358 \$1235 \$1132 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$360 \$1236 \$1131 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$362 \$1236 \$1134 \$1035 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$364 \$1235 \$1135 \$1035 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P
+ PS=10.82U PD=10.82U
M$366 vdd \$1134 \$1135 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$367 vdd \$1025 \$1136 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$368 \$1136 \$1023 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$369 vdd \$1021 \$1137 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$370 \$1137 \$1019 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$371 \$1237 \$1137 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$373 \$1237 \$1136 \$866 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$375 vdd \$1035 \$1138 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$376 \$1138 \$787 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$377 fout \$1138 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$378 \$1238 fout \$790 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$380 \$1238 define vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$382 \$1624 \$1442 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$383 \$1442 fin vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$384 \$1904 \$473 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$385 \$1444 \$1442 \$1443 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$386 \$1443 \$1624 \$1904 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$387 vdd \$1508 \$1444 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$388 \$1508 \$1443 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$389 \$1444 \$1445 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$390 \$1446 \$1442 \$1508 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$391 vdd vss \$1445 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$392 vdd \$1446 \$1509 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$393 \$1447 \$1624 \$1446 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$394 vdd \$1509 \$1447 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$395 \$1509 \$1445 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$396 \$1448 \$1509 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$397 vdd \$1905 \$1513 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$398 vdd \$473 \$1905 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$399 \$1449 \$1448 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$401 \$1449 \$738 \$1450 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$403 \$1905 \$1451 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$404 \$1451 \$1450 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$405 vdd \$473 \$1906 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$406 vdd \$1510 \$473 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$407 \$1907 \$473 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$408 \$1511 \$1636 \$1907 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$409 \$473 \$1511 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$410 \$1510 vss vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$411 \$1452 \$1363 \$1511 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$412 vdd \$1510 \$1908 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$413 vdd \$1512 \$1452 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$414 \$1453 \$1636 \$1512 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$415 \$1908 \$1452 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$416 \$1512 \$1363 \$1908 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$417 vdd \$1513 \$1453 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$418 vdd fin \$1363 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$419 vdd \$1363 \$1636 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$420 \$1625 \$1454 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$421 \$1454 \$473 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$422 \$1909 \$1515 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$423 \$1456 \$1454 \$1455 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$424 vdd \$1514 \$1456 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$425 \$1455 \$1625 \$1909 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$426 \$1514 \$1455 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$427 \$1456 \$1457 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$428 \$1458 \$1454 \$1514 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$429 vdd \$1 \$1457 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$430 vdd \$1458 \$1515 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$431 \$1459 \$1625 \$1458 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$432 vdd \$1515 \$1459 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$433 \$1515 \$1457 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$434 \$1091 pd1 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$435 \$1094 \$1515 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$436 \$1626 \$1460 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$437 \$1460 \$1094 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$438 \$1910 \$1517 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$439 \$1462 \$1460 \$1461 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$440 \$1461 \$1626 \$1910 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$441 vdd \$1516 \$1462 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$442 \$1516 \$1461 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$443 \$1462 \$1463 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$444 \$1464 \$1460 \$1516 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$445 vdd \$1 \$1463 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$446 vdd \$1464 \$1517 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$447 \$1465 \$1626 \$1464 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$448 vdd \$1517 \$1465 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$449 \$1517 \$1463 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$450 \$1099 \$1517 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$451 \$1096 pd2 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$452 \$1627 \$1466 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$453 \$1466 \$1099 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$454 \$1911 \$1519 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$455 \$1468 \$1466 \$1467 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$456 \$1467 \$1627 \$1911 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$457 vdd \$1518 \$1468 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$458 \$1518 \$1467 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$459 \$1468 \$1469 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$460 \$1470 \$1466 \$1518 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$461 vdd \$1 \$1469 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$462 vdd \$1470 \$1519 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$463 \$1471 \$1627 \$1470 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$464 vdd \$1519 \$1471 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$465 \$1519 \$1469 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$466 \$1104 \$1519 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$467 \$1101 pd3 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$468 \$1628 \$1472 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$469 \$1472 \$1104 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$470 \$1912 \$1521 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$471 \$1474 \$1472 \$1473 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$472 \$1473 \$1628 \$1912 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$473 vdd \$1520 \$1474 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$474 \$1520 \$1473 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$475 \$1474 \$1475 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$476 \$1476 \$1472 \$1520 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$477 vdd \$1 \$1475 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$478 vdd \$1476 \$1521 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$479 \$1477 \$1628 \$1476 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$480 vdd \$1521 \$1477 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$481 \$1521 \$1475 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$482 \$1106 pd4 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$483 \$1109 \$1521 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$484 \$1629 \$1478 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$485 \$1478 \$1109 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$486 \$1913 \$1523 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$487 \$1480 \$1478 \$1479 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$488 vdd \$1522 \$1480 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$489 \$1479 \$1629 \$1913 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$490 \$1522 \$1479 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$491 \$1480 \$1481 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$492 \$1482 \$1478 \$1522 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$493 vdd \$1 \$1481 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$494 vdd \$1482 \$1523 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$495 \$1483 \$1629 \$1482 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$496 vdd \$1523 \$1483 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$497 \$1523 \$1481 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$498 \$1114 \$1523 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$499 \$1111 pd5 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$500 \$1630 \$1484 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$501 \$1484 \$1114 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$502 \$1914 \$1525 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$503 \$1486 \$1484 \$1485 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$504 vdd \$1524 \$1486 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$505 \$1485 \$1630 \$1914 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$506 \$1524 \$1485 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$507 \$1486 \$1487 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$508 \$1488 \$1484 \$1524 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$509 vdd \$1 \$1487 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$510 vdd \$1488 \$1525 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$511 \$1489 \$1630 \$1488 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$512 vdd \$1525 \$1489 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$513 \$1525 \$1487 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$514 \$1116 pd6 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$515 \$1119 \$1525 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$516 \$1631 \$1490 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$517 \$1490 \$1119 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$518 \$1915 \$1527 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$519 \$1492 \$1490 \$1491 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$520 vdd \$1526 \$1492 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$521 \$1491 \$1631 \$1915 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$522 \$1526 \$1491 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$523 \$1492 \$1493 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$524 \$1494 \$1490 \$1526 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$525 vdd \$1 \$1493 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$526 vdd \$1494 \$1527 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$527 \$1495 \$1631 \$1494 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$528 vdd \$1527 \$1495 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$529 \$1527 \$1493 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$530 \$1121 pd7 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$531 \$1124 \$1527 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$532 \$1632 \$1496 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$533 \$1496 \$1124 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$534 \$1916 \$1529 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$535 \$1498 \$1496 \$1497 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$536 vdd \$1528 \$1498 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$537 \$1497 \$1632 \$1916 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$538 \$1528 \$1497 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$539 \$1498 \$1499 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$540 \$1500 \$1496 \$1528 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$541 vdd \$1 \$1499 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$542 vdd \$1500 \$1529 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$543 \$1501 \$1632 \$1500 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$544 vdd \$1529 \$1501 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$545 \$1529 \$1499 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$546 \$1129 \$1529 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$547 \$1126 pd8 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$548 \$1633 \$1502 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$549 \$1502 \$1129 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$550 \$1917 \$1531 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$551 \$1504 \$1502 \$1503 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$552 vdd \$1530 \$1504 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$553 \$1503 \$1633 \$1917 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$554 \$1530 \$1503 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$555 \$1504 \$1505 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$556 \$1506 \$1502 \$1530 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$557 vdd \$1 \$1505 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$558 vdd \$1506 \$1531 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$559 \$1507 \$1633 \$1506 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$560 vdd \$1531 \$1507 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$561 \$1531 \$1505 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$562 \$1134 \$1531 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$563 \$1131 pd9 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$564 vss sd9 \$77 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$565 \$226 \$119 \$78 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$567 \$226 \$120 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$569 \$79 \$80 \$120 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$570 vss \$121 \$79 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$571 \$81 \$3 \$121 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$572 vss \$78 \$81 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$573 vss \$3 \$80 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$574 vss sd8 \$4 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$575 \$227 \$123 \$82 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$577 \$227 \$124 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$579 \$83 \$84 \$124 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$580 vss \$125 \$83 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$581 \$85 \$5 \$125 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$582 vss \$82 \$85 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$583 vss \$5 \$84 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$584 vss sd7 \$86 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$585 \$228 \$127 \$87 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$587 \$228 \$128 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$589 \$88 \$89 \$128 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$590 vss \$129 \$88 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$591 \$90 \$6 \$129 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$592 vss \$87 \$90 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$593 vss \$6 \$89 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$594 vss sd6 \$91 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$595 \$229 \$454 \$131 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$597 \$229 \$132 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$599 \$92 \$93 \$132 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$600 vss \$133 \$92 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$601 \$94 \$7 \$133 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$602 vss \$131 \$94 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$603 vss \$7 \$93 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$604 vss sd5 \$8 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$605 \$230 \$458 \$135 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$607 \$230 \$136 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$609 \$95 \$96 \$136 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$610 vss \$137 \$95 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$611 \$97 \$9 \$137 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$612 vss \$135 \$97 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$613 vss \$9 \$96 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$614 vss sd4 \$98 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$615 \$231 \$139 \$99 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$617 \$231 \$140 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$619 \$100 \$101 \$140 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$620 vss \$141 \$100 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$621 \$102 \$10 \$141 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$622 vss \$99 \$102 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$623 vss \$10 \$101 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$624 vss sd3 \$103 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$625 \$232 \$143 \$104 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$627 \$232 \$144 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$629 \$105 \$106 \$144 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$630 vss \$145 \$105 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$631 \$107 \$11 \$145 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$632 vss \$104 \$107 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$633 vss \$11 \$106 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$634 vss sd2 \$108 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$635 \$233 \$468 \$109 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$637 \$233 \$147 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$639 \$110 \$111 \$147 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$640 vss \$148 \$110 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$641 \$112 \$12 \$148 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$642 vss \$109 \$112 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$643 vss \$12 \$111 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$644 vss sd1 \$113 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$645 \$234 \$150 \$114 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$647 \$234 \$151 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$649 \$115 \$116 \$151 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$650 vss \$152 \$115 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$651 \$117 \$13 \$152 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$652 vss \$114 \$117 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$653 vss \$13 \$116 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$654 vss \$78 \$443 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$655 \$444 \$78 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$656 \$120 \$3 \$444 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$657 \$119 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$658 \$371 \$119 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$660 \$371 \$79 \$445 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$662 \$121 \$80 \$445 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$663 vss \$446 \$3 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$664 vss \$82 \$446 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$665 \$447 \$82 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$666 \$124 \$5 \$447 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$667 \$123 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$668 \$372 \$123 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$670 \$372 \$83 \$448 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$672 \$125 \$84 \$448 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$673 vss \$449 \$5 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$674 vss \$87 \$449 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$675 \$450 \$87 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$676 \$128 \$6 \$450 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$677 \$127 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$678 \$373 \$127 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$680 \$373 \$88 \$451 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$682 \$129 \$89 \$451 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$683 vss \$452 \$6 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$684 vss \$131 \$452 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$685 \$453 \$131 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$686 \$132 \$7 \$453 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$687 \$454 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$688 \$374 \$454 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$690 \$374 \$92 \$455 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$692 \$133 \$93 \$455 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$693 vss \$456 \$7 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$694 vss \$135 \$456 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$695 \$457 \$135 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$696 \$136 \$9 \$457 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$697 \$458 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$698 \$375 \$458 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$700 \$375 \$95 \$459 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$702 \$137 \$96 \$459 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$703 vss \$460 \$9 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$704 vss \$99 \$460 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$705 \$461 \$99 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$706 \$140 \$10 \$461 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$707 \$139 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$708 \$376 \$139 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$710 \$376 \$100 \$462 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$712 \$141 \$101 \$462 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$713 vss \$463 \$10 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$714 vss \$104 \$463 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$715 \$464 \$104 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$716 \$144 \$11 \$464 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$717 \$143 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$718 \$377 \$143 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$720 \$377 \$105 \$465 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$722 \$145 \$106 \$465 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$723 vss \$466 \$11 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$724 vss \$109 \$466 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$725 \$467 \$109 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$726 \$147 \$12 \$467 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$727 \$468 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$728 \$378 \$468 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$730 \$378 \$110 \$469 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$732 \$148 \$111 \$469 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$733 vss \$470 \$12 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$734 vss \$114 \$470 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$735 \$471 \$114 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$736 \$151 \$13 \$471 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$737 \$150 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$738 \$379 \$150 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$740 \$379 \$115 \$472 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$742 \$152 \$116 \$472 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$743 vss \$473 \$13 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$744 vss \$788 \$738 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$745 \$738 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$746 vss \$741 \$740 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$747 \$868 \$789 \$741 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$749 \$868 \$681 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$751 vss \$745 \$742 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$752 \$742 \$744 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$753 \$869 \$689 \$744 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$755 \$869 \$688 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$757 \$870 \$687 \$745 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$759 \$870 \$686 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$761 \$746 \$443 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$762 \$871 \$746 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$764 \$872 \$443 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$766 \$871 \$77 \$681 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$768 \$872 \$749 \$681 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$770 vss \$77 \$749 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$771 \$750 \$446 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$772 \$873 \$750 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$774 \$874 \$446 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$776 \$873 \$4 \$682 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$778 \$874 \$753 \$682 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$780 vss \$4 \$753 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$781 \$754 \$449 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$782 \$875 \$754 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$784 \$876 \$449 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$786 \$875 \$86 \$683 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$788 \$876 \$757 \$683 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$790 vss \$86 \$757 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$791 \$758 \$452 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$792 \$877 \$758 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$794 \$878 \$452 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$796 \$877 \$91 \$684 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$798 \$878 \$761 \$684 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$800 vss \$91 \$761 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$801 \$762 \$456 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$802 \$879 \$762 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$804 \$880 \$456 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$806 \$879 \$8 \$685 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$808 \$880 \$765 \$685 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$810 vss \$8 \$765 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$811 \$766 \$460 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$812 \$881 \$766 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$814 \$882 \$460 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$816 \$881 \$98 \$686 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$818 \$882 \$769 \$686 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$820 vss \$98 \$769 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$821 \$770 \$463 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$822 \$883 \$770 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$824 \$884 \$463 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$826 \$883 \$103 \$687 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$828 \$884 \$773 \$687 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$830 vss \$103 \$773 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$831 \$774 \$466 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$832 \$885 \$774 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$834 \$886 \$466 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$836 \$885 \$108 \$688 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$838 \$886 \$777 \$688 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$840 vss \$108 \$777 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$841 \$778 \$470 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$842 \$887 \$778 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$844 \$888 \$470 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$846 \$887 \$113 \$689 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$848 \$888 \$781 \$689 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$850 vss \$113 \$781 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$851 \$889 \$1033 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$853 \$889 \$1031 \$782 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$855 \$890 \$1029 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$857 \$890 \$1027 \$783 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$859 vss \$783 \$785 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$860 \$785 \$782 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$861 \$891 \$785 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$863 \$891 \$866 \$786 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$865 \$787 \$786 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$866 vss \$790 \$1 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$867 vss \$740 \$788 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$868 \$788 \$738 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$869 vss \$1088 \$789 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$870 \$1015 \$742 \$1088 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$872 \$1015 \$1089 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$874 vss \$1016 \$1089 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$875 \$1089 \$1090 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$876 \$1017 \$685 \$1090 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$878 \$1017 \$684 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$880 \$1018 \$683 \$1016 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$882 \$1018 \$682 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$884 \$1092 \$1091 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$885 \$1020 \$1092 \$1019 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$887 \$1093 \$1091 \$1019 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$889 \$1020 \$1094 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$891 \$1093 \$1095 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$893 vss \$1094 \$1095 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$894 \$1097 \$1096 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$895 \$1022 \$1097 \$1021 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$897 \$1098 \$1096 \$1021 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$899 \$1022 \$1099 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$901 \$1098 \$1100 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$903 vss \$1099 \$1100 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$904 \$1102 \$1101 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$905 \$1024 \$1102 \$1023 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$907 \$1103 \$1101 \$1023 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$909 \$1024 \$1104 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$911 \$1103 \$1105 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$913 vss \$1104 \$1105 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$914 \$1107 \$1106 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$915 \$1026 \$1107 \$1025 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$917 \$1108 \$1106 \$1025 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$919 \$1026 \$1109 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$921 \$1108 \$1110 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$923 vss \$1109 \$1110 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$924 \$1112 \$1111 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$925 \$1028 \$1112 \$1027 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$927 \$1113 \$1111 \$1027 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$929 \$1028 \$1114 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$931 \$1113 \$1115 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$933 vss \$1114 \$1115 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$934 \$1117 \$1116 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$935 \$1030 \$1117 \$1029 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$937 \$1118 \$1116 \$1029 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$939 \$1030 \$1119 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$941 \$1118 \$1120 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$943 vss \$1119 \$1120 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$944 \$1122 \$1121 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$945 \$1032 \$1122 \$1031 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$947 \$1123 \$1121 \$1031 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$949 \$1032 \$1124 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$951 \$1123 \$1125 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$953 vss \$1124 \$1125 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$954 \$1127 \$1126 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$955 \$1034 \$1127 \$1033 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$957 \$1128 \$1126 \$1033 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$959 \$1034 \$1129 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$961 \$1128 \$1130 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$963 vss \$1129 \$1130 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$964 \$1132 \$1131 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$965 \$1036 \$1132 \$1035 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$967 \$1133 \$1131 \$1035 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$969 \$1036 \$1134 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$971 \$1133 \$1135 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$973 vss \$1134 \$1135 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$974 \$1037 \$1025 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$976 \$1037 \$1023 \$1136 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$978 \$1038 \$1021 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$980 \$1038 \$1019 \$1137 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$982 vss \$1137 \$866 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$983 \$866 \$1136 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$984 \$1039 \$1035 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$986 \$1039 \$787 \$1138 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$988 fout \$1138 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$989 vss fout \$790 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$990 \$790 define vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$991 \$1624 \$1442 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$992 \$1442 fin vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$993 \$1904 \$473 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$994 \$1444 \$1624 \$1443 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$995 \$1443 \$1442 \$1904 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$996 \$1634 \$1508 \$1444 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$998 \$1508 \$1443 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$999 \$1634 \$1445 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1001 \$1446 \$1624 \$1508 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1002 vss vss \$1445 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1003 \$1892 \$1446 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1005 \$1447 \$1442 \$1446 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1006 \$1892 \$1445 \$1509 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1008 vss \$1509 \$1447 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1009 \$1448 \$1509 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1010 vss \$1905 \$1513 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1011 \$1893 \$473 \$1905 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1013 vss \$1448 \$1450 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1014 \$1893 \$1451 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1016 \$1450 \$738 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1017 \$1451 \$1450 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1018 vss \$473 \$1906 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1019 \$1635 \$1510 \$473 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1021 \$1907 \$473 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1022 \$1511 \$1363 \$1907 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1023 \$1635 \$1511 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1025 \$1510 vss vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1026 \$1452 \$1636 \$1511 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1027 \$1894 \$1510 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1029 vss \$1512 \$1452 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1030 \$1894 \$1452 \$1908 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1032 \$1453 \$1363 \$1512 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1033 \$1512 \$1636 \$1908 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1034 vss \$1513 \$1453 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1035 vss fin \$1363 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1036 vss \$1363 \$1636 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1037 \$1625 \$1454 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1038 \$1454 \$473 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1039 \$1909 \$1515 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1040 \$1456 \$1625 \$1455 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1041 \$1455 \$1454 \$1909 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1042 \$1637 \$1514 \$1456 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1044 \$1514 \$1455 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1045 \$1637 \$1457 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1047 \$1458 \$1625 \$1514 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1048 vss \$1 \$1457 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1049 \$1895 \$1458 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1051 \$1459 \$1454 \$1458 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1052 \$1895 \$1457 \$1515 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1054 vss \$1515 \$1459 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1055 \$1094 \$1515 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1056 \$1091 pd1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1057 \$1626 \$1460 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1058 \$1460 \$1094 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1059 \$1910 \$1517 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1060 \$1462 \$1626 \$1461 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1061 \$1638 \$1516 \$1462 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1063 \$1461 \$1460 \$1910 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1064 \$1516 \$1461 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1065 \$1638 \$1463 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1067 \$1464 \$1626 \$1516 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1068 vss \$1 \$1463 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1069 \$1896 \$1464 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1071 \$1465 \$1460 \$1464 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1072 \$1896 \$1463 \$1517 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1074 vss \$1517 \$1465 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1075 \$1099 \$1517 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1076 \$1096 pd2 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1077 \$1627 \$1466 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1078 \$1466 \$1099 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1079 \$1911 \$1519 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1080 \$1468 \$1627 \$1467 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1081 \$1467 \$1466 \$1911 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1082 \$1639 \$1518 \$1468 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1084 \$1518 \$1467 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1085 \$1639 \$1469 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1087 \$1470 \$1627 \$1518 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1088 vss \$1 \$1469 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1089 \$1897 \$1470 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1091 \$1471 \$1466 \$1470 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1092 \$1897 \$1469 \$1519 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1094 vss \$1519 \$1471 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1095 \$1104 \$1519 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1096 \$1101 pd3 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1097 \$1628 \$1472 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1098 \$1472 \$1104 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1099 \$1912 \$1521 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1100 \$1474 \$1628 \$1473 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1101 \$1473 \$1472 \$1912 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1102 \$1640 \$1520 \$1474 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1104 \$1520 \$1473 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1105 \$1640 \$1475 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1107 \$1476 \$1628 \$1520 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1108 vss \$1 \$1475 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1109 \$1898 \$1476 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1111 \$1477 \$1472 \$1476 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1112 \$1898 \$1475 \$1521 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1114 vss \$1521 \$1477 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1115 \$1109 \$1521 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1116 \$1106 pd4 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1117 \$1629 \$1478 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1118 \$1478 \$1109 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1119 \$1913 \$1523 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1120 \$1480 \$1629 \$1479 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1121 \$1641 \$1522 \$1480 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1123 \$1479 \$1478 \$1913 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1124 \$1522 \$1479 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1125 \$1641 \$1481 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1127 \$1482 \$1629 \$1522 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1128 vss \$1 \$1481 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1129 \$1899 \$1482 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1131 \$1483 \$1478 \$1482 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1132 \$1899 \$1481 \$1523 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1134 vss \$1523 \$1483 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1135 \$1114 \$1523 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1136 \$1111 pd5 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1137 \$1630 \$1484 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1138 \$1484 \$1114 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1139 \$1914 \$1525 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1140 \$1486 \$1630 \$1485 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1141 \$1485 \$1484 \$1914 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1142 \$1642 \$1524 \$1486 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1144 \$1524 \$1485 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1145 \$1642 \$1487 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1147 \$1488 \$1630 \$1524 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1148 vss \$1 \$1487 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1149 \$1900 \$1488 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1151 \$1489 \$1484 \$1488 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1152 \$1900 \$1487 \$1525 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1154 vss \$1525 \$1489 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1155 \$1119 \$1525 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1156 \$1116 pd6 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1157 \$1631 \$1490 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1158 \$1490 \$1119 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1159 \$1915 \$1527 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1160 \$1492 \$1631 \$1491 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1161 \$1643 \$1526 \$1492 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1163 \$1491 \$1490 \$1915 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1164 \$1526 \$1491 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1165 \$1643 \$1493 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1167 \$1494 \$1631 \$1526 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1168 vss \$1 \$1493 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1169 \$1901 \$1494 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1171 \$1495 \$1490 \$1494 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1172 \$1901 \$1493 \$1527 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1174 vss \$1527 \$1495 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1175 \$1124 \$1527 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1176 \$1121 pd7 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1177 \$1632 \$1496 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1178 \$1496 \$1124 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1179 \$1916 \$1529 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1180 \$1498 \$1632 \$1497 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1181 \$1644 \$1528 \$1498 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1183 \$1497 \$1496 \$1916 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1184 \$1528 \$1497 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1185 \$1644 \$1499 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1187 \$1500 \$1632 \$1528 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1188 vss \$1 \$1499 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1189 \$1902 \$1500 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1191 \$1501 \$1496 \$1500 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1192 \$1902 \$1499 \$1529 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1194 vss \$1529 \$1501 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1195 \$1126 pd8 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1196 \$1129 \$1529 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1197 \$1633 \$1502 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1198 \$1502 \$1129 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1199 \$1917 \$1531 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1200 \$1504 \$1633 \$1503 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1201 \$1645 \$1530 \$1504 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1203 \$1503 \$1502 \$1917 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1204 \$1530 \$1503 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1205 \$1645 \$1505 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1207 \$1506 \$1633 \$1530 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1208 vss \$1 \$1505 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1209 \$1903 \$1506 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$1211 \$1507 \$1502 \$1506 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$1212 \$1903 \$1505 \$1531 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P
+ PS=4.74U PD=4.74U
M$1214 vss \$1531 \$1507 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1215 \$1131 pd9 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$1216 \$1134 \$1531 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
.ENDS asc_dual_psd_def_20250809
