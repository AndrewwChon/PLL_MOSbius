** sch_path: /foss/designs/libs/xp_core_analog/asc_PFD_DFF/asc_PFD_DFF.sch
.subckt asc_PFD_DFF vdd vss down up fref fdiv
*.PININFO vdd:B vss:B fref:B fdiv:B up:B down:B
x1 fref vdd net3 vdd vss up rst asc_dff_rst
x2 fdiv vdd net4 vdd vss down rst asc_dff_rst
x4 net2 vdd net1 vss inv1u05u
x3 net1 vss rst vdd asc_delay
x5 vdd net2 up down vss asc_NAND
.ends

* expanding   symbol:  libs/core_analog/asc_dff_rst/asc_dff_rst.sym # of pins=7
** sym_path: /foss/designs/libs/core_analog/asc_dff_rst/asc_dff_rst.sym
** sch_path: /foss/designs/libs/core_analog/asc_dff_rst/asc_dff_rst.sch
.subckt asc_dff_rst clk D Qb vdd vss Q rst
*.PININFO clk:B vdd:B vss:B D:B Q:B Qb:B rst:B
x1 net3 vdd net2 vss inv1u05u
x2 clk vdd clkb vss inv1u05u
x3 net1 vss clkb net3 clka vdd pass1u05u
x5 net3 vss clka net6 clkb vdd pass1u05u
x6 net2 vss clka net5 clkb vdd pass1u05u
x8 Qb vdd net4 vss inv1u05u
x9 net5 vss clkb net4 clka vdd pass1u05u
x10 clkb vdd clka vss inv1u05u
x11 D vdd net1 vss inv1u05u
x12 Qb vdd Q vss inv1u05u
x13 rst vdd rstb vss inv1u05u
x4 vdd net6 net2 rstb vss asc_NAND
x7 vdd Qb rstb net5 vss asc_NAND
.ends


* expanding   symbol:  libs/core_analog/inv1u05u/inv1u05u.sym # of pins=4
** sym_path: /foss/designs/libs/core_analog/inv1u05u/inv1u05u.sym
** sch_path: /foss/designs/libs/core_analog/inv1u05u/inv1u05u.sch
.subckt inv1u05u in vdd out vss
*.PININFO in:B out:B vss:B vdd:B
M1 out in vdd vdd pfet_03v3 L=0.5u W=3.0u nf=1 m=1
M2 out in vss vss nfet_03v3 L=0.5u W=1.0u nf=1 m=1
.ends


* expanding   symbol:  libs/core_analog/asc_delay/asc_delay.sym # of pins=4
** sym_path: /foss/designs/libs/core_analog/asc_delay/asc_delay.sym
** sch_path: /foss/designs/libs/core_analog/asc_delay/asc_delay.sch
.subckt asc_delay in vss out vdd
*.PININFO vdd:B vss:B in:B out:B
x1 in vdd net1 vss inv1u05u
x2 net1 vdd out vss inv1u05u
.ends


* expanding   symbol:  libs/core_analog/asc_NAND/asc_NAND.sym # of pins=5
** sym_path: /foss/designs/libs/core_analog/asc_NAND/asc_NAND.sym
** sch_path: /foss/designs/libs/core_analog/asc_NAND/asc_NAND.sch
.subckt asc_NAND VDD OUT A B VSS
*.PININFO VDD:B VSS:B B:B A:B OUT:B
M1 OUT A net1 VSS nfet_03v3 L=0.5u W=2u nf=1 m=1
M2 OUT A VDD VDD pfet_03v3 L=0.5u W=3u nf=1 m=1
M3 net1 B VSS VSS nfet_03v3 L=0.5u W=2u nf=1 m=1
M4 OUT B VDD VDD pfet_03v3 L=0.5u W=3u nf=1 m=1
.ends


* expanding   symbol:  libs/core_analog/pass1u05u/pass1u05u.sym # of pins=6
** sym_path: /foss/designs/libs/core_analog/pass1u05u/pass1u05u.sym
** sch_path: /foss/designs/libs/core_analog/pass1u05u/pass1u05u.sch
.subckt pass1u05u ind vss clkn ins clkp vdd
*.PININFO ind:B ins:B clkn:B clkp:B vdd:B vss:B
M1 ind clkp ins vdd pfet_03v3 L=0.5u W=3.0u nf=1 m=1
M2 ind clkn ins vss nfet_03v3 L=0.5u W=1.0u nf=1 m=1
.ends

