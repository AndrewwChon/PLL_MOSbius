* NGSPICE file created from SRegister_10.ext - technology: gf180mcuD

.subckt gf180mcu_fd_sc_mcu9t5v0__and2_1 A1 A2 VDD VSS Z VNW VPW
X0 VDD A2 a_36_201# VNW pfet_05v0 ad=0.5054p pd=2.57u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1 a_244_201# A1 a_36_201# VPW nfet_05v0 ad=0.1056p pd=0.98u as=0.2904p ps=2.2u w=0.66u l=0.6u
X2 Z a_36_201# VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.3894p ps=2.06u w=1.32u l=0.6u
X3 Z a_36_201# VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.5054p ps=2.57u w=1.83u l=0.5u
X4 VSS A2 a_244_201# VPW nfet_05v0 ad=0.3894p pd=2.06u as=0.1056p ps=0.98u w=0.66u l=0.6u
X5 a_36_201# A1 VDD VNW pfet_05v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__latq_1$1 D E Q VDD VSS VNW VPW
X0 VSS a_1020_652# Q VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X1 a_504_110# a_36_92# VDD VNW pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X2 VDD a_1020_652# Q VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X3 a_1264_107# a_36_92# a_1020_652# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X4 VSS E a_36_92# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X5 VSS a_1364_532# a_1264_107# VPW nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X6 VDD E a_36_92# VNW pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X7 VDD a_1364_532# a_1224_652# VNW pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X8 a_872_652# D VDD VNW pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X9 a_1364_532# a_1020_652# VDD VNW pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X10 a_1020_652# a_504_110# a_872_107# VPW nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X11 a_872_107# D VSS VPW nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X12 a_1020_652# a_36_92# a_872_652# VNW pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X13 a_504_110# a_36_92# VSS VPW nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X14 a_1364_532# a_1020_652# VSS VPW nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X15 a_1224_652# a_504_110# a_1020_652# VNW pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt DFF_2phase_1 D Q PHI_1 PHI_2 VSSd VDDd
Xgf180mcu_fd_sc_mcu9t5v0__latq_1$1_0 gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1/Q PHI_2 Q
+ VDDd VSSd VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1$1
Xgf180mcu_fd_sc_mcu9t5v0__latq_1$1_1 D PHI_1 gf180mcu_fd_sc_mcu9t5v0__latq_1$1_1/Q
+ VDDd VSSd VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1$1
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1 I VDD VSS ZN VNW VPW
X0 ZN I VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__or2_1 A1 A2 VDD VSS Z VNW VPW
X0 a_255_756# A1 a_67_756# VNW pfet_05v0 ad=0.2379p pd=1.435u as=0.4026p ps=2.71u w=0.915u l=0.5u
X1 VSS A2 a_67_756# VPW nfet_05v0 ad=0.3828p pd=2.08u as=0.1716p ps=1.18u w=0.66u l=0.6u
X2 VDD A2 a_255_756# VNW pfet_05v0 ad=0.57645p pd=2.69u as=0.2379p ps=1.435u w=0.915u l=0.5u
X3 Z a_67_756# VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.3828p ps=2.08u w=1.32u l=0.6u
X4 Z a_67_756# VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.57645p ps=2.69u w=1.83u l=0.5u
X5 a_67_756# A1 VSS VPW nfet_05v0 ad=0.1716p pd=1.18u as=0.2904p ps=2.2u w=0.66u l=0.6u
.ends

.subckt Register_unitcell out d en default phi2 phi1 q VDDd VSSd
Xgf180mcu_fd_sc_mcu9t5v0__and2_1_1 q en VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1_0/A2
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1
XDFF_2phase_1_0 d q phi1 phi2 VSSd VDDd DFF_2phase_1
Xgf180mcu_fd_sc_mcu9t5v0__inv_1_0 en VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1_0/ZN
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1
Xgf180mcu_fd_sc_mcu9t5v0__or2_1_0 gf180mcu_fd_sc_mcu9t5v0__or2_1_0/A1 gf180mcu_fd_sc_mcu9t5v0__or2_1_0/A2
+ VDDd VSSd out VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1
Xgf180mcu_fd_sc_mcu9t5v0__and2_1_0 gf180mcu_fd_sc_mcu9t5v0__inv_1_0/ZN default VDDd
+ VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1_0/A1 VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1
.ends

.subckt SRegister_10 VDDd VSSd out[1] out[2] out[3] out[4] out[5] out[6] out[7] out[8]
+ out[9] out[10] d q default10 default9 default8 default7 default6 default5 default4
+ default3 default2 default1 phi1 phi2 en
XRegister_unitcell_0 out[2] Register_unitcell_6/q en default2 phi2 phi1 Register_unitcell_7/d
+ VDDd VSSd Register_unitcell
XRegister_unitcell_1 out[6] Register_unitcell_9/q en default6 phi2 phi1 Register_unitcell_2/d
+ VDDd VSSd Register_unitcell
XRegister_unitcell_2 out[7] Register_unitcell_2/d en default7 phi2 phi1 Register_unitcell_3/d
+ VDDd VSSd Register_unitcell
XRegister_unitcell_3 out[8] Register_unitcell_3/d en default8 phi2 phi1 Register_unitcell_4/d
+ VDDd VSSd Register_unitcell
XRegister_unitcell_5 out[10] Register_unitcell_5/d en default10 phi2 phi1 q VDDd VSSd
+ Register_unitcell
XRegister_unitcell_4 out[9] Register_unitcell_4/d en default9 phi2 phi1 Register_unitcell_5/d
+ VDDd VSSd Register_unitcell
XRegister_unitcell_6 out[1] d en default1 phi2 phi1 Register_unitcell_6/q VDDd VSSd
+ Register_unitcell
XRegister_unitcell_7 out[3] Register_unitcell_7/d en default3 phi2 phi1 Register_unitcell_8/d
+ VDDd VSSd Register_unitcell
XRegister_unitcell_8 out[4] Register_unitcell_8/d en default4 phi2 phi1 Register_unitcell_9/d
+ VDDd VSSd Register_unitcell
XRegister_unitcell_9 out[5] Register_unitcell_9/d en default5 phi2 phi1 Register_unitcell_9/q
+ VDDd VSSd Register_unitcell
.ends

