* NGSPICE file created from top_level_nosc_20250831.ext - technology: gf180mcuD

.subckt nfet$47 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$46 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$50 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$49 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$48 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$47 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$51 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$50 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$49 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$48 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt asc_drive_buffer_up vss vdd out in
Xnfet$47_0 m1_778_712# vss m1_506_712# m1_506_712# m1_506_712# m1_778_712# m1_778_712#
+ vss m1_506_712# vss nfet$47
Xpfet$46_0 out out m1_778_712# vdd m1_778_712# out vdd vdd m1_778_712# out m1_778_712#
+ m1_778_712# out m1_778_712# vdd m1_778_712# vdd m1_778_712# pfet$46
Xnfet$50_0 m1_n566_1318# vss m1_n30_1318# vss nfet$50
Xpfet$49_0 vdd vdd m1_n30_1318# m1_n566_1318# pfet$49
Xnfet$48_0 out out vss m1_778_712# m1_778_712# out vss m1_778_712# m1_778_712# m1_778_712#
+ out m1_778_712# m1_778_712# out vss m1_778_712# vss vss nfet$48
Xpfet$47_0 m1_778_712# vdd vdd m1_778_712# m1_506_712# m1_506_712# m1_778_712# vdd
+ m1_506_712# m1_506_712# pfet$47
Xnfet$51_0 in vss m1_n566_1318# vss nfet$51
Xpfet$50_0 vdd vdd m1_n566_1318# in pfet$50
Xnfet$49_0 m1_n30_1318# vss m1_506_712# vss nfet$49
Xpfet$48_0 vdd vdd m1_506_712# m1_n30_1318# pfet$48
.ends

.subckt nfet$79 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$93 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$87 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$86 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$68 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$66 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$78 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$91 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$103 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$71 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$77 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$74 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$84 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$90 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$100 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$83 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$101 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$76 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$69 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$82 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$75 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$81 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$74 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$78 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$98 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$80 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$67 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$94 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$97 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$77 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$108 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$72 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$96 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$89 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$95 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$88 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$106 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$70 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$87 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$93 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$86 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$104 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$92 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$79 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$85 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$91 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$81 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$76 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$84 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$102 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$90 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$83 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$82 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$75 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$99 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$80 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$109 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$73 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$97 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$96 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$89 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$107 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$95 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$88 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$94 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$105 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$92 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$85 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt asc_dual_psd_def_20250809 vdd vss pd1 pd2 pd3 pd4 pd5 pd6 pd7 pd8 pd9 fout
+ sd1 sd2 sd3 sd4 sd5 sd6 sd7 sd8 sd9 fin define w_n11156_26804#
Xnfet$79_1 m1_n3218_15478# vss m1_4620_20152# vss nfet$79
Xnfet$93_3 m1_11381_15778# m1_11381_15778# m1_11271_18030# m1_11271_18030# m1_11507_17358#
+ vss nfet$93
Xpfet$87_4 w_n11156_26804# m1_n2567_23922# m1_n3184_24224# m1_n4464_25980# pfet$87
Xnfet$86_2 m1_8154_21786# m1_8154_21786# vss vss m1_6992_21586# vss nfet$86
Xpfet$68_25 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_17526_19550# m1_13514_15478#
+ m1_13514_15478# pfet$68
Xpfet$68_14 w_n11156_26804# m1_n927_19404# m1_n927_19404# m1_n59_19550# m1_n7383_17599#
+ m1_n7383_17599# pfet$68
Xpfet$66_9 w_n11156_26804# w_n11156_26804# m1_8172_15778# m1_5302_17714# pfet$66
Xpfet$78_0 w_n11156_26804# m1_34093_22102# w_n11156_26804# m1_28490_22513# pfet$78
Xnfet$91_0 m1_34093_22102# vss fout vss nfet$91
Xpfet_0 w_n11156_26804# w_n11156_26804# m1_3049_25662# m1_2912_25858# pfet
Xnfet$103_1 m1_n10796_25662# m1_n10572_23922# m1_n10308_24542# vss nfet$103
Xpfet$71_7 w_n11156_26804# w_n11156_26804# m1_11654_20152# m1_5148_15478# pfet$71
Xnfet$93_26 m1_14127_16080# m1_14127_16080# m1_13668_17714# m1_13668_17714# m1_14225_16398#
+ vss nfet$93
Xnfet$77_49 m1_21564_17714# vss m1_18665_17343# vss nfet$77
Xnfet$77_27 m1_1119_17714# vss m1_3989_15778# vss nfet$77
Xnfet$77_16 m1_6275_17836# m1_7198_15778# m1_6377_16202# vss nfet$77
Xnfet$77_38 m1_n2250_17343# m1_n1989_16202# m1_n2474_17518# vss nfet$77
Xnfet$93_15 m1_n1989_16202# m1_n1989_16202# vss vss m1_n2507_16398# vss nfet$93
Xpfet_91 w_n11156_26804# w_n11156_26804# m1_23356_21786# pd8 pfet
Xpfet_80 w_n11156_26804# w_n11156_26804# m1_17058_24346# m1_n7513_20152# pfet
Xnfet$74_39 pd4 vss m1_9288_21786# vss nfet$74
Xpfet$66_91 w_n11156_26804# m1_24287_16080# m1_23820_18030# m1_22848_17343# pfet$66
Xpfet$66_80 w_n11156_26804# w_n11156_26804# m1_15564_15778# m1_15921_16080# pfet$66
Xnfet$74_28 m1_3394_25858# vss m1_4005_21786# vss nfet$74
Xnfet$74_17 m1_11639_23922# vss m1_12259_24224# vss nfet$74
Xnfet$93_4 m1_10560_16202# m1_10560_16202# vss vss m1_10042_16398# vss nfet$93
Xpfet$87_5 w_n11156_26804# m1_n10572_23922# m1_n10308_24542# m1_n10933_25858# pfet$87
Xnfet$86_3 m1_7522_21786# m1_7522_21786# vss vss m1_6360_21586# vss nfet$86
Xnfet$79_2 m1_n7401_15478# vss m1_1103_20152# vss nfet$79
Xpfet$68_26 w_n11156_26804# m1_n1927_20274# m1_n1927_20274# m1_17526_19550# m1_13198_17714#
+ m1_13198_17714# pfet$68
Xpfet$68_15 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_n59_19550# m1_n7401_15478#
+ m1_n7401_15478# pfet$68
Xpfet$78_1 w_n11156_26804# w_n11156_26804# m1_34093_22102# m1_34843_21786# pfet$78
Xnfet$84_0 pd1 vss m1_n1263_21786# vss nfet$84
Xnfet$103_2 m1_n10933_25858# m1_n10309_25662# m1_n10572_23922# vss nfet$103
Xpfet_1 w_n11156_26804# m1_3536_25662# m1_3273_23922# m1_3049_25662# pfet
Xpfet$90_0 w_n11156_26804# w_n11156_26804# m1_n8145_21908# m1_n6839_20152# pfet$90
Xpfet$71_8 w_n11156_26804# w_n11156_26804# m1_n1133_19550# m1_n7383_17599# pfet$71
Xnfet$93_27 m1_18310_16080# m1_18310_16080# vss vss m1_19873_17358# vss nfet$93
Xnfet$93_16 m1_19747_15778# m1_19747_15778# m1_19637_18030# m1_19637_18030# m1_19873_17358#
+ vss nfet$93
Xnfet$77_28 m1_1933_17343# vss m1_2092_17836# vss nfet$77
Xnfet$77_17 m1_649_17714# vss m1_n2250_17343# vss nfet$77
Xnfet$77_39 m1_n3064_17714# vss m1_n3534_17714# vss nfet$77
Xpfet_92 w_n11156_26804# w_n11156_26804# m1_28492_25858# m1_29607_24346# pfet
Xpfet_81 w_n11156_26804# w_n11156_26804# m1_18339_24542# m1_15943_25858# pfet
Xpfet_70 w_n11156_26804# w_n11156_26804# m1_14156_24542# m1_11760_25858# pfet
Xnfet$74_29 m1_15943_25858# vss m1_14556_21786# vss nfet$74
Xpfet$66_92 w_n11156_26804# m1_15454_18030# w_n11156_26804# m1_14127_16080# pfet$66
Xpfet$66_81 w_n11156_26804# w_n11156_26804# m1_13668_17714# m1_14127_16080# pfet$66
Xpfet$66_70 w_n11156_26804# w_n11156_26804# m1_18824_17836# m1_18665_17343# pfet$66
Xnfet$74_18 m1_7095_25858# vss m1_7232_25662# vss nfet$74
Xnfet$100_10 m1_9624_19404# m1_9624_19404# vss vss m1_n3724_21430# vss nfet$100
Xpfet$87_6 w_n11156_26804# m1_n8848_25658# m1_n8055_24542# m1_n10796_25662# pfet$87
Xnfet$79_3 m1_649_17714# vss m1_5901_19550# vss nfet$79
Xnfet$93_5 m1_9944_16080# m1_9944_16080# m1_9485_17714# m1_9485_17714# m1_10042_16398#
+ vss nfet$93
Xnfet$86_4 m1_1120_21786# m1_1120_21786# vss vss m1_n42_21586# vss nfet$86
Xpfet$68_27 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_20407_19850# m1_22205_20152#
+ m1_22205_20152# pfet$68
Xpfet$68_16 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_28077_19550# m1_26063_15478#
+ m1_26063_15478# pfet$68
Xpfet$78_2 w_n11156_26804# w_n11156_26804# m1_30256_22102# m1_7388_22513# pfet$78
Xnfet$84_1 pd2 vss m1_2254_21786# vss nfet$84
Xnfet$77_0 m1_9485_17714# vss m1_9015_17714# vss nfet$77
Xnfet$103_3 m1_n10796_25662# m1_n9952_24224# m1_n8848_25658# vss nfet$103
Xpfet$71_9 w_n11156_26804# w_n11156_26804# m1_27003_19550# m1_25747_17714# pfet$71
Xpfet_2 w_n11156_26804# w_n11156_26804# m1_3394_25858# m1_4509_24346# pfet
Xnfet$93_17 m1_22493_16080# m1_22493_16080# vss vss m1_24056_17358# vss nfet$93
Xnfet$77_29 m1_3372_16080# vss m1_3015_15778# vss nfet$77
Xnfet$77_18 m1_1119_17714# vss m1_649_17714# vss nfet$77
Xpfet$83_0 w_n11156_26804# w_n11156_26804# m1_n7247_17714# m1_n6788_16080# pfet$83
Xpfet$90_1 w_n11156_26804# m1_n5227_20152# w_n11156_26804# m1_n1927_20274# pfet$90
Xnfet$101_0 m1_n8625_26174# vss m1_n8055_24542# vss nfet$101
Xpfet_93 w_n11156_26804# m1_28991_24224# m1_30095_25658# m1_28010_25858# pfet
Xpfet_82 w_n11156_26804# w_n11156_26804# m1_21241_24346# m1_n7513_20152# pfet
Xpfet_71 w_n11156_26804# w_n11156_26804# m1_11039_21786# m1_11760_25858# pfet
Xpfet_60 w_n11156_26804# w_n11156_26804# m1_20126_25858# m1_21241_24346# pfet
Xpfet$66_93 w_n11156_26804# m1_23820_18030# w_n11156_26804# m1_22493_16080# pfet$66
Xpfet$66_82 w_n11156_26804# m1_13668_17714# w_n11156_26804# m1_14743_16202# pfet$66
Xpfet$66_71 w_n11156_26804# w_n11156_26804# m1_19747_15778# m1_20104_16080# pfet$66
Xpfet$66_60 w_n11156_26804# w_n11156_26804# m1_n194_15778# m1_n3064_17714# pfet$66
Xnfet$74_19 m1_7456_23922# vss m1_8076_24224# vss nfet$74
Xnfet$100_11 m1_n6380_21786# m1_n6380_21786# m1_n6839_21786# m1_n6839_21786# m1_n6282_21430#
+ vss nfet$100
Xnfet$79_4 m1_4832_17714# vss m1_9418_19550# vss nfet$79
Xnfet$93_6 m1_1578_16080# m1_1578_16080# vss vss m1_3141_17358# vss nfet$93
Xpfet$87_7 w_n11156_26804# m1_n3541_23922# m1_n4362_24346# m1_n4623_25487# pfet$87
Xnfet$86_5 m1_4005_21786# m1_4005_21786# vss vss m1_2843_21586# vss nfet$86
Xpfet$68_28 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_21043_19550# m1_17697_15478#
+ m1_17697_15478# pfet$68
Xpfet$68_17 w_n11156_26804# m1_n3822_20130# m1_n3822_20130# m1_28077_19550# m1_25747_17714#
+ m1_25747_17714# pfet$68
Xpfet$78_3 w_n11156_26804# m1_31535_22102# w_n11156_26804# m1_3871_22513# pfet$78
Xnfet$84_2 pd9 vss m1_26873_21786# vss nfet$84
Xnfet$77_1 m1_9015_17714# vss m1_6116_17343# vss nfet$77
Xnfet$103_4 m1_n4623_25487# m1_n2567_23922# m1_n3184_24224# vss nfet$103
Xpfet_3 w_n11156_26804# m1_3394_25858# w_n11156_26804# m1_4997_25658# pfet
Xnfet$93_18 m1_23930_15778# m1_23930_15778# m1_23820_18030# m1_23820_18030# m1_24056_17358#
+ vss nfet$93
Xpfet$76_0 w_n11156_26804# m1_32818_20470# m1_32818_20470# m1_33050_19550# m1_30256_19792#
+ m1_30256_19792# pfet$76
Xnfet$77_19 m1_n7513_20152# vss m1_1578_16080# vss nfet$77
Xpfet$90_2 w_n11156_26804# w_n11156_26804# m1_n5227_20152# m1_n2543_20130# pfet$90
Xpfet$83_1 w_n11156_26804# m1_n7247_17714# w_n11156_26804# m1_n6172_16202# pfet$83
Xnfet$101_1 m1_n8625_26174# vss m1_n7082_23622# vss nfet$101
Xpfet_94 w_n11156_26804# m1_28492_25858# w_n11156_26804# m1_30095_25658# pfet
Xpfet_83 w_n11156_26804# m1_21729_25658# m1_22522_24542# m1_19781_25662# pfet
Xpfet_72 w_n11156_26804# m1_13363_25658# m1_14156_24542# m1_11415_25662# pfet
Xpfet_61 w_n11156_26804# m1_24452_24542# w_n11156_26804# m1_25424_24346# pfet
Xpfet_50 w_n11156_26804# w_n11156_26804# m1_20268_25662# m1_20126_25858# pfet
Xpfet$66_50 w_n11156_26804# m1_n1168_15778# m1_n1989_16202# m1_n2250_17343# pfet$66
Xpfet$66_94 w_n11156_26804# w_n11156_26804# m1_22624_17518# m1_22034_17714# pfet$66
Xpfet$66_83 w_n11156_26804# m1_16538_15778# m1_15921_16080# m1_14641_17836# pfet$66
Xpfet$66_72 w_n11156_26804# m1_20721_15778# m1_20104_16080# m1_18824_17836# pfet$66
Xpfet$66_61 w_n11156_26804# m1_n811_16080# m1_n1278_18030# m1_n2250_17343# pfet$66
Xnfet$79_5 m1_965_15478# vss m1_8137_20152# vss nfet$79
Xnfet$93_7 m1_5761_16080# m1_5761_16080# m1_5302_17714# m1_5302_17714# m1_5859_16398#
+ vss nfet$93
Xnfet$86_6 m1_4637_21786# m1_4637_21786# vss vss m1_3475_21586# vss nfet$86
Xpfet$68_29 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_23924_19850# m1_25722_20152#
+ m1_25722_20152# pfet$68
Xpfet$68_18 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_27441_19850# m1_29239_20152#
+ m1_29239_20152# pfet$68
Xpfet$78_4 w_n11156_26804# m1_30256_22102# w_n11156_26804# m1_9645_21447# pfet$78
Xnfet$77_2 m1_6275_17836# m1_7555_16080# m1_7088_18030# vss nfet$77
Xnfet$103_5 m1_n4464_25980# m1_n3541_23922# m1_n4362_24346# vss nfet$103
Xpfet_4 w_n11156_26804# w_n11156_26804# m1_3893_24224# m1_3273_23922# pfet
Xpfet$76_1 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_33050_19550# m1_31535_19792#
+ m1_31535_19792# pfet$76
Xpfet$90_3 w_n11156_26804# m1_n4485_20152# w_n11156_26804# m1_n3206_20274# pfet$90
Xpfet$83_2 w_n11156_26804# w_n11156_26804# m1_n5461_18030# m1_n5351_15778# pfet$83
Xpfet$69_0 w_n11156_26804# w_n11156_26804# m1_n1133_21590# m1_n1263_21786# pfet$69
Xnfet$82_0 m1_n10452_25858# vss m1_n1271_25858# vss nfet$82
Xnfet$93_19 m1_23109_16202# m1_23109_16202# vss vss m1_22591_16398# vss nfet$93
Xnfet$101_2 vss vss m1_n9336_24346# vss nfet$101
Xpfet_95 w_n11156_26804# w_n11156_26804# m1_28991_24224# m1_28371_23922# pfet
Xpfet_84 w_n11156_26804# w_n11156_26804# m1_23827_25858# m1_18073_21786# pfet
Xpfet_73 w_n11156_26804# m1_16086_24542# w_n11156_26804# m1_17058_24346# pfet
Xpfet_62 w_n11156_26804# w_n11156_26804# m1_24452_24542# m1_24808_24224# pfet
Xpfet_51 w_n11156_26804# w_n11156_26804# m1_20625_24224# m1_20005_23922# pfet
Xpfet_40 w_n11156_26804# w_n11156_26804# m1_11760_25858# m1_12875_24346# pfet
Xpfet$66_95 w_n11156_26804# w_n11156_26804# m1_21564_17714# m1_22034_17714# pfet$66
Xpfet$66_84 w_n11156_26804# w_n11156_26804# m1_17381_17714# m1_17851_17714# pfet$66
Xpfet$66_73 w_n11156_26804# w_n11156_26804# m1_16538_15778# m1_13668_17714# pfet$66
Xpfet$66_62 w_n11156_26804# w_n11156_26804# m1_23007_17836# m1_22848_17343# pfet$66
Xpfet$66_40 w_n11156_26804# m1_10560_16202# m1_10075_17518# m1_10458_17836# pfet$66
Xpfet$66_51 w_n11156_26804# w_n11156_26804# m1_n1168_15778# m1_n811_16080# pfet$66
Xnfet$86_7 m1_488_21786# m1_488_21786# vss vss m1_n674_21586# vss nfet$86
Xnfet$79_6 m1_9015_17714# vss m1_12935_19550# vss nfet$79
Xnfet$93_8 m1_3015_15778# m1_3015_15778# m1_2905_18030# m1_2905_18030# m1_3141_17358#
+ vss nfet$93
Xpfet$68_19 w_n11156_26804# m1_n3822_20130# m1_n3822_20130# m1_27441_19850# m1_27003_19550#
+ m1_27003_19550# pfet$68
Xpfet$78_5 w_n11156_26804# w_n11156_26804# m1_31535_22102# m1_354_22513# pfet$78
Xnfet$77_3 m1_n7513_20152# vss m1_9944_16080# vss nfet$77
Xpfet_5 w_n11156_26804# m1_3893_24224# m1_4997_25658# m1_2912_25858# pfet
Xnfet$103_6 m1_n4464_25980# m1_n3184_24224# m1_n3651_26174# vss nfet$103
Xpfet$76_2 w_n11156_26804# m1_32818_21586# m1_32818_21586# m1_33050_22344# m1_30256_22102#
+ m1_30256_22102# pfet$76
Xpfet$90_4 w_n11156_26804# m1_n6839_20152# w_n11156_26804# m1_n927_19404# pfet$90
Xpfet$83_3 w_n11156_26804# m1_n5461_18030# w_n11156_26804# m1_n6788_16080# pfet$83
Xnfet$75_0 m1_n1133_21590# m1_n1133_21590# m1_354_22513# m1_354_22513# m1_n674_21586#
+ vss nfet$75
Xnfet$101_3 fin vss m1_n10933_25858# vss nfet$101
Xnfet$82_1 m1_n789_25858# vss m1_n647_25662# vss nfet$82
Xpfet$69_1 w_n11156_26804# w_n11156_26804# m1_11671_21786# m1_11039_21786# pfet$69
Xpfet_110 w_n11156_26804# m1_11903_24542# w_n11156_26804# m1_12875_24346# pfet
Xpfet_96 w_n11156_26804# m1_28635_24542# w_n11156_26804# m1_29607_24346# pfet
Xpfet$81_0 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_36073_22344# define
+ define pfet$81
Xpfet_85 w_n11156_26804# m1_24188_23922# m1_24452_24542# m1_23827_25858# pfet
Xpfet_74 w_n11156_26804# w_n11156_26804# m1_14556_21786# m1_15943_25858# pfet
Xpfet_63 w_n11156_26804# w_n11156_26804# m1_19781_25662# m1_19644_25858# pfet
Xpfet_52 w_n11156_26804# m1_20268_25662# m1_20005_23922# m1_19781_25662# pfet
Xpfet_41 w_n11156_26804# w_n11156_26804# m1_9288_21786# pd4 pfet
Xpfet_30 w_n11156_26804# w_n11156_26804# m1_2912_25858# m1_488_21786# pfet
Xpfet$66_96 w_n11156_26804# w_n11156_26804# m1_18665_17343# m1_21564_17714# pfet$66
Xpfet$66_85 w_n11156_26804# m1_18926_16202# m1_18441_17518# m1_18824_17836# pfet$66
Xpfet$66_74 w_n11156_26804# w_n11156_26804# m1_14641_17836# m1_14482_17343# pfet$66
Xpfet$66_63 w_n11156_26804# m1_23930_15778# m1_23109_16202# m1_22848_17343# pfet$66
Xpfet$66_30 w_n11156_26804# w_n11156_26804# m1_1933_17343# m1_4832_17714# pfet$66
Xpfet$66_41 w_n11156_26804# w_n11156_26804# m1_10075_17518# m1_9485_17714# pfet$66
Xpfet$66_52 w_n11156_26804# m1_n3064_17714# w_n11156_26804# m1_n1989_16202# pfet$66
Xnfet$75_10 m1_19839_21786# m1_19839_21786# m1_21456_22513# m1_21456_22513# m1_21060_21586#
+ vss nfet$75
Xnfet$86_8 m1_25739_21786# m1_25739_21786# vss vss m1_24577_21586# vss nfet$86
Xnfet$93_9 m1_2194_16202# m1_2194_16202# vss vss m1_1676_16398# vss nfet$93
Xnfet$79_7 m1_5148_15478# vss m1_11654_20152# vss nfet$79
Xpfet$66_110 w_n11156_26804# w_n11156_26804# m1_10458_17836# m1_10299_17343# pfet$66
Xnfet$77_4 m1_10299_17343# m1_10560_16202# m1_10075_17518# vss nfet$77
Xnfet$103_7 m1_n4623_25487# m1_n4362_24346# m1_n4847_25662# vss nfet$103
Xpfet_6 w_n11156_26804# w_n11156_26804# m1_3536_25662# m1_3394_25858# pfet
Xpfet$90_5 w_n11156_26804# w_n11156_26804# m1_n4485_20152# m1_n3822_20130# pfet$90
Xpfet$76_3 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_33050_22344# m1_31535_22102#
+ m1_31535_22102# pfet$76
Xpfet$83_4 w_n11156_26804# w_n11156_26804# m1_26217_17714# m1_26676_16080# pfet$83
Xnfet$75_1 m1_n1263_21786# m1_n1263_21786# m1_354_22513# m1_354_22513# m1_n42_21586#
+ vss nfet$75
Xnfet$82_2 m1_n1271_25858# vss m1_n1134_25662# vss nfet$82
Xpfet$69_2 w_n11156_26804# w_n11156_26804# m1_12935_21590# m1_12805_21786# pfet$69
Xnfet$101_4 m1_n10572_23922# vss m1_n9952_24224# vss nfet$101
Xpfet_100 w_n11156_26804# w_n11156_26804# m1_29607_24346# m1_n7513_20152# pfet
Xpfet_97 w_n11156_26804# w_n11156_26804# m1_21590_21786# m1_24309_25858# pfet
Xpfet_86 w_n11156_26804# m1_28634_25662# m1_28371_23922# m1_28147_25662# pfet
Xpfet$81_1 w_n11156_26804# m1_35837_22102# m1_35837_22102# m1_36073_22344# fout fout
+ pfet$81
Xpfet_75 w_n11156_26804# w_n11156_26804# m1_19644_25858# m1_14556_21786# pfet
Xpfet_64 w_n11156_26804# w_n11156_26804# m1_22522_24542# m1_20126_25858# pfet
Xpfet_53 w_n11156_26804# m1_20625_24224# m1_21729_25658# m1_19644_25858# pfet
Xpfet_42 w_n11156_26804# m1_11760_25858# w_n11156_26804# m1_13363_25658# pfet
Xpfet_31 w_n11156_26804# m1_3273_23922# m1_3537_24542# m1_2912_25858# pfet
Xpfet_20 w_n11156_26804# w_n11156_26804# m1_4509_24346# m1_n7513_20152# pfet
Xpfet$74_0 w_n11156_26804# w_n11156_26804# m1_n646_24542# m1_n290_24224# pfet$74
Xnfet$78_10 m1_21590_21786# vss m1_22222_21786# vss nfet$78
Xpfet$66_97 w_n11156_26804# w_n11156_26804# m1_22493_16080# m1_n7513_20152# pfet$66
Xpfet$66_86 w_n11156_26804# m1_19637_18030# w_n11156_26804# m1_18310_16080# pfet$66
Xpfet$66_75 w_n11156_26804# w_n11156_26804# m1_17697_15478# sd3 pfet$66
Xpfet$66_64 w_n11156_26804# w_n11156_26804# m1_23930_15778# m1_24287_16080# pfet$66
Xpfet$66_20 w_n11156_26804# w_n11156_26804# m1_1119_17714# m1_1578_16080# pfet$66
Xpfet$66_31 w_n11156_26804# m1_3372_16080# m1_2905_18030# m1_1933_17343# pfet$66
Xpfet$66_42 w_n11156_26804# m1_11271_18030# w_n11156_26804# m1_9944_16080# pfet$66
Xpfet$66_53 w_n11156_26804# w_n11156_26804# m1_n3218_15478# sd8 pfet$66
Xnfet$75_11 m1_19969_21590# m1_19969_21590# m1_21456_22513# m1_21456_22513# m1_20428_21586#
+ vss nfet$75
Xnfet$86_9 m1_25107_21786# m1_25107_21786# vss vss m1_23945_21586# vss nfet$86
Xnfet$79_8 m1_n7383_17599# vss m1_n1133_19550# vss nfet$79
Xnfet$98_0 m1_n10452_25858# m1_n10452_25858# m1_n7186_25858# m1_n7186_25858# m1_n6629_25502#
+ vss nfet$98
Xnfet$86_10 m1_21590_21786# m1_21590_21786# vss vss m1_20428_21586# vss nfet$86
Xpfet$66_100 w_n11156_26804# w_n11156_26804# m1_23820_18030# m1_23930_15778# pfet$66
Xnfet$77_5 m1_10458_17836# m1_11738_16080# m1_11271_18030# vss nfet$77
Xpfet_7 w_n11156_26804# w_n11156_26804# m1_7232_25662# m1_7095_25858# pfet
Xpfet$83_5 w_n11156_26804# m1_26217_17714# w_n11156_26804# m1_27292_16202# pfet$83
Xnfet$82_3 m1_n7513_20152# vss m1_326_24346# vss nfet$82
Xpfet$90_6 w_n11156_26804# w_n11156_26804# m1_n6839_20152# m1_n6973_21481# pfet$90
Xnfet$75_2 m1_9288_21786# m1_9288_21786# m1_9645_21447# m1_9645_21447# m1_10509_21586#
+ vss nfet$75
Xpfet$69_3 w_n11156_26804# w_n11156_26804# m1_9418_21590# m1_9288_21786# pfet$69
Xnfet$101_5 m1_n10933_25858# vss m1_n10796_25662# vss nfet$101
Xpfet_65 w_n11156_26804# w_n11156_26804# m1_18073_21786# m1_20126_25858# pfet
Xpfet_54 w_n11156_26804# w_n11156_26804# m1_24808_24224# m1_24188_23922# pfet
Xpfet_43 w_n11156_26804# w_n11156_26804# m1_12805_21786# pd5 pfet
Xpfet$71_10 w_n11156_26804# w_n11156_26804# m1_29239_20152# m1_26063_15478# pfet$71
Xpfet_32 w_n11156_26804# w_n11156_26804# m1_7720_24542# m1_8076_24224# pfet
Xpfet_21 w_n11156_26804# m1_7456_23922# m1_7720_24542# m1_7095_25858# pfet
Xpfet_10 w_n11156_26804# m1_8076_24224# m1_9180_25658# m1_7095_25858# pfet
Xpfet$74_1 w_n11156_26804# m1_n789_25858# w_n11156_26804# m1_814_25658# pfet$74
Xpfet_101 w_n11156_26804# w_n11156_26804# m1_28010_25858# m1_21590_21786# pfet
Xpfet_98 w_n11156_26804# m1_30095_25658# m1_30888_24542# m1_28147_25662# pfet
Xpfet_87 w_n11156_26804# w_n11156_26804# m1_28147_25662# m1_28010_25858# pfet
Xpfet_76 w_n11156_26804# m1_20005_23922# m1_20269_24542# m1_19644_25858# pfet
Xnfet$78_11 m1_18073_21786# vss m1_18705_21786# vss nfet$78
Xnfet$80_0 sd9 vss m1_n7401_15478# vss nfet$80
Xpfet$67_0 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_n674_22102# m1_n1133_21590#
+ m1_n1133_21590# pfet$67
Xpfet$66_98 w_n11156_26804# m1_20104_16080# m1_19637_18030# m1_18665_17343# pfet$66
Xpfet$66_87 w_n11156_26804# w_n11156_26804# m1_18310_16080# m1_n7513_20152# pfet$66
Xnfet$94_10 m1_9331_15478# m1_9331_15478# m1_n3822_21786# m1_n3822_21786# m1_13373_20470#
+ vss nfet$94
Xpfet$66_76 w_n11156_26804# m1_17851_17714# w_n11156_26804# m1_18926_16202# pfet$66
Xpfet$66_65 w_n11156_26804# m1_24904_15778# m1_24287_16080# m1_23007_17836# pfet$66
Xpfet$66_21 w_n11156_26804# w_n11156_26804# m1_965_15478# sd7 pfet$66
Xpfet$66_10 w_n11156_26804# m1_8172_15778# m1_7555_16080# m1_6275_17836# pfet$66
Xpfet$66_32 w_n11156_26804# w_n11156_26804# m1_2905_18030# m1_3015_15778# pfet$66
Xpfet$66_43 w_n11156_26804# w_n11156_26804# m1_11271_18030# m1_11381_15778# pfet$66
Xpfet$66_54 w_n11156_26804# w_n11156_26804# m1_n1278_18030# m1_n1168_15778# pfet$66
Xnfet$75_12 m1_16322_21786# m1_16322_21786# m1_17939_22513# m1_17939_22513# m1_17543_21586#
+ vss nfet$75
Xnfet$79_9 m1_25747_17714# vss m1_27003_19550# vss nfet$79
Xpfet$66_101 w_n11156_26804# w_n11156_26804# m1_19637_18030# m1_19747_15778# pfet$66
Xnfet$98_1 m1_n6111_25858# m1_n6111_25858# vss vss m1_n6629_25502# vss nfet$98
Xnfet$86_11 m1_22222_21786# m1_22222_21786# vss vss m1_21060_21586# vss nfet$86
Xnfet$77_6 m1_6116_17343# vss m1_6275_17836# vss nfet$77
Xpfet$97_0 w_n11156_26804# w_n11156_26804# m1_n8145_21908# m1_n6839_20152# pfet$97
Xpfet_8 w_n11156_26804# w_n11156_26804# m1_8076_24224# m1_7456_23922# pfet
Xpfet$69_10 w_n11156_26804# w_n11156_26804# m1_23486_21590# m1_23356_21786# pfet$69
Xpfet$83_6 w_n11156_26804# w_n11156_26804# m1_28003_18030# m1_28113_15778# pfet$83
Xnfet$82_4 m1_n789_25858# vss m1_1607_24542# vss nfet$82
Xpfet$90_7 w_n11156_26804# m1_n6839_21786# w_n11156_26804# m1_n5764_21786# pfet$90
Xnfet$75_3 m1_9418_21590# m1_9418_21590# m1_9645_21447# m1_9645_21447# m1_9877_21586#
+ vss nfet$75
Xpfet$69_4 w_n11156_26804# w_n11156_26804# m1_8154_21786# m1_7522_21786# pfet$69
Xnfet$101_6 m1_n10452_25858# vss m1_n10309_25662# vss nfet$101
Xpfet$71_11 w_n11156_26804# w_n11156_26804# m1_18688_20152# m1_13514_15478# pfet$71
Xpfet_102 w_n11156_26804# m1_28371_23922# m1_28635_24542# m1_28010_25858# pfet
Xpfet_99 w_n11156_26804# w_n11156_26804# m1_26705_24542# m1_24309_25858# pfet
Xpfet_88 w_n11156_26804# w_n11156_26804# m1_28634_25662# m1_28492_25858# pfet
Xpfet_77 w_n11156_26804# w_n11156_26804# m1_20269_24542# m1_20625_24224# pfet
Xpfet_66 w_n11156_26804# w_n11156_26804# m1_15461_25858# m1_11039_21786# pfet
Xpfet_55 w_n11156_26804# m1_24451_25662# m1_24188_23922# m1_23964_25662# pfet
Xpfet_44 w_n11156_26804# m1_15943_25858# w_n11156_26804# m1_17546_25658# pfet
Xnfet$80_1 sd2 vss m1_21880_15478# vss nfet$80
Xpfet_33 w_n11156_26804# w_n11156_26804# m1_7522_21786# m1_7577_25858# pfet
Xpfet_22 w_n11156_26804# w_n11156_26804# m1_3537_24542# m1_3893_24224# pfet
Xpfet_11 w_n11156_26804# w_n11156_26804# m1_7719_25662# m1_7577_25858# pfet
Xpfet$74_2 w_n11156_26804# w_n11156_26804# m1_n789_25858# m1_326_24346# pfet$74
Xpfet$67_1 w_n11156_26804# m1_7388_22513# m1_7388_22513# m1_6988_22402# m1_7522_21786#
+ m1_7522_21786# pfet$67
Xnfet$78_12 m1_14556_21786# vss m1_15188_21786# vss nfet$78
Xnfet$94_11 m1_15171_20152# m1_15171_20152# m1_n3822_21786# m1_n3822_21786# m1_14005_20470#
+ vss nfet$94
Xpfet$66_22 w_n11156_26804# w_n11156_26804# m1_3015_15778# m1_3372_16080# pfet$66
Xpfet$66_11 w_n11156_26804# w_n11156_26804# m1_9485_17714# m1_9944_16080# pfet$66
Xpfet$66_33 w_n11156_26804# w_n11156_26804# m1_5892_17518# m1_5302_17714# pfet$66
Xpfet$66_44 w_n11156_26804# w_n11156_26804# m1_649_17714# m1_1119_17714# pfet$66
Xpfet$66_55 w_n11156_26804# w_n11156_26804# m1_n2474_17518# m1_n3064_17714# pfet$66
Xpfet$66_99 w_n11156_26804# m1_23109_16202# m1_22624_17518# m1_23007_17836# pfet$66
Xpfet$66_88 w_n11156_26804# w_n11156_26804# m1_18441_17518# m1_17851_17714# pfet$66
Xpfet$66_77 w_n11156_26804# w_n11156_26804# m1_17851_17714# m1_18310_16080# pfet$66
Xpfet$66_66 w_n11156_26804# w_n11156_26804# m1_24904_15778# m1_22034_17714# pfet$66
Xpfet$77_10 w_n11156_26804# m1_30256_22102# w_n11156_26804# m1_9645_21447# pfet$77
Xnfet$75_13 m1_16452_21590# m1_16452_21590# m1_17939_22513# m1_17939_22513# m1_16911_21586#
+ vss nfet$75
Xpfet$66_102 w_n11156_26804# w_n11156_26804# m1_13198_17714# m1_13668_17714# pfet$66
Xnfet_20 m1_21241_24346# m1_21241_24346# m1_20126_25858# m1_20126_25858# m1_22188_25502#
+ vss nfet
Xnfet$86_12 m1_18073_21786# m1_18073_21786# vss vss m1_16911_21586# vss nfet$86
Xnfet$77_7 m1_9485_17714# vss m1_10075_17518# vss nfet$77
Xpfet$90_10 w_n11156_26804# w_n11156_26804# m1_n5227_21418# m1_6107_19404# pfet$90
Xpfet_9 w_n11156_26804# m1_7719_25662# m1_7456_23922# m1_7232_25662# pfet
Xnfet$108_0 m1_n5227_20152# vss m1_n6380_21786# vss nfet$108
Xpfet$69_11 w_n11156_26804# w_n11156_26804# m1_18705_21786# m1_18073_21786# pfet$69
Xpfet$83_7 w_n11156_26804# m1_28003_18030# w_n11156_26804# m1_26676_16080# pfet$83
Xnfet$82_5 m1_n789_25858# vss m1_488_21786# vss nfet$82
Xpfet$90_8 w_n11156_26804# m1_n4485_21904# w_n11156_26804# m1_9624_19404# pfet$90
Xpfet$69_5 w_n11156_26804# w_n11156_26804# m1_1120_21786# m1_488_21786# pfet$69
Xnfet$75_4 m1_5901_21590# m1_5901_21590# m1_7388_22513# m1_7388_22513# m1_6360_21586#
+ vss nfet$75
Xnfet$101_7 m1_n7320_25516# vss m1_n2567_23922# vss nfet$101
Xpfet$71_12 w_n11156_26804# w_n11156_26804# m1_15171_20152# m1_9331_15478# pfet$71
Xnfet$80_2 sd1 vss m1_26063_15478# vss nfet$80
Xpfet_103 w_n11156_26804# w_n11156_26804# m1_28635_24542# m1_28991_24224# pfet
Xpfet_89 w_n11156_26804# w_n11156_26804# m1_19839_21786# pd7 pfet
Xpfet_78 w_n11156_26804# m1_20269_24542# w_n11156_26804# m1_21241_24346# pfet
Xpfet_67 w_n11156_26804# m1_15822_23922# m1_16086_24542# m1_15461_25858# pfet
Xpfet_56 w_n11156_26804# m1_24808_24224# m1_25912_25658# m1_23827_25858# pfet
Xpfet_45 w_n11156_26804# w_n11156_26804# m1_16442_24224# m1_15822_23922# pfet
Xpfet$74_3 w_n11156_26804# m1_n646_24542# w_n11156_26804# m1_326_24346# pfet$74
Xpfet_34 w_n11156_26804# m1_9180_25658# m1_9973_24542# m1_7232_25662# pfet
Xpfet_23 w_n11156_26804# m1_3537_24542# w_n11156_26804# m1_4509_24346# pfet
Xpfet_12 w_n11156_26804# m1_7577_25858# w_n11156_26804# m1_9180_25658# pfet
Xpfet$67_2 w_n11156_26804# m1_7388_22513# m1_7388_22513# m1_6360_22102# m1_8154_21786#
+ m1_8154_21786# pfet$67
Xnfet$78_13 m1_16322_21786# vss m1_16452_21590# vss nfet$78
Xnfet$94_12 m1_18688_20152# m1_18688_20152# m1_n1927_20274# m1_n1927_20274# m1_17522_20470#
+ vss nfet$94
Xpfet$66_89 w_n11156_26804# w_n11156_26804# m1_22848_17343# m1_25747_17714# pfet$66
Xpfet$66_78 w_n11156_26804# w_n11156_26804# m1_13514_15478# sd4 pfet$66
Xpfet$66_67 w_n11156_26804# m1_22034_17714# w_n11156_26804# m1_23109_16202# pfet$66
Xpfet$66_12 w_n11156_26804# m1_3989_15778# m1_3372_16080# m1_2092_17836# pfet$66
Xpfet$66_23 w_n11156_26804# m1_5302_17714# w_n11156_26804# m1_6377_16202# pfet$66
Xpfet$66_34 w_n11156_26804# w_n11156_26804# m1_5761_16080# m1_n7513_20152# pfet$66
Xpfet$66_45 w_n11156_26804# w_n11156_26804# m1_9944_16080# m1_n7513_20152# pfet$66
Xpfet$66_56 w_n11156_26804# m1_n1278_18030# w_n11156_26804# m1_n2605_16080# pfet$66
Xpfet$72_0 w_n11156_26804# w_n11156_26804# m1_n7401_15478# sd9 pfet$72
Xpfet$77_11 w_n11156_26804# w_n11156_26804# m1_30256_22102# m1_7388_22513# pfet$77
Xnfet$75_14 m1_12805_21786# m1_12805_21786# m1_14422_22513# m1_14422_22513# m1_14026_21586#
+ vss nfet$75
Xnfet_21 m1_28991_24224# m1_28991_24224# m1_28635_24542# m1_28635_24542# m1_29089_24542#
+ vss nfet
Xnfet_10 m1_17546_25658# m1_17546_25658# vss vss m1_18005_25502# vss nfet
Xnfet$86_13 m1_18705_21786# m1_18705_21786# vss vss m1_17543_21586# vss nfet$86
Xpfet$66_103 w_n11156_26804# m1_14743_16202# m1_14258_17518# m1_14641_17836# pfet$66
Xnfet$77_8 m1_7555_16080# vss m1_7198_15778# vss nfet$77
Xpfet$90_11 w_n11156_26804# w_n11156_26804# m1_n4485_21904# m1_n3822_21786# pfet$90
Xnfet$96_0 m1_n6274_17836# m1_n4994_16080# m1_n5461_18030# vss nfet$96
Xpfet$69_12 w_n11156_26804# w_n11156_26804# m1_16452_21590# m1_16322_21786# pfet$69
Xnfet$108_1 m1_n4485_20152# m1_n6380_21786# vss vss nfet$108
Xpfet$90_9 w_n11156_26804# m1_n5227_21418# w_n11156_26804# m1_2590_19404# pfet$90
Xpfet$69_6 w_n11156_26804# w_n11156_26804# m1_5901_21590# m1_5771_21786# pfet$69
Xnfet$82_6 m1_n910_23922# vss m1_n290_24224# vss nfet$82
Xnfet$75_5 m1_2254_21786# m1_2254_21786# m1_3871_22513# m1_3871_22513# m1_3475_21586#
+ vss nfet$75
Xnfet$101_8 m1_n4623_25487# vss m1_n4464_25980# vss nfet$101
Xpfet$71_13 w_n11156_26804# w_n11156_26804# m1_16452_19550# m1_13198_17714# pfet$71
Xpfet_104 w_n11156_26804# m1_25912_25658# m1_26705_24542# m1_23964_25662# pfet
Xpfet$74_4 w_n11156_26804# w_n11156_26804# m1_32675_25947# m1_33790_24346# pfet$74
Xpfet_79 w_n11156_26804# m1_17546_25658# m1_18339_24542# m1_15598_25662# pfet
Xpfet_68 w_n11156_26804# w_n11156_26804# m1_16086_24542# m1_16442_24224# pfet
Xpfet_57 w_n11156_26804# w_n11156_26804# m1_24451_25662# m1_24309_25858# pfet
Xpfet_46 w_n11156_26804# m1_16442_24224# m1_17546_25658# m1_15461_25858# pfet
Xpfet_35 w_n11156_26804# m1_7720_24542# w_n11156_26804# m1_8692_24346# pfet
Xpfet_24 w_n11156_26804# w_n11156_26804# m1_5790_24542# m1_3394_25858# pfet
Xpfet_13 w_n11156_26804# w_n11156_26804# m1_12259_24224# m1_11639_23922# pfet
Xpfet$67_3 w_n11156_26804# m1_9645_21447# m1_9645_21447# m1_10505_22402# m1_11039_21786#
+ m1_11039_21786# pfet$67
Xnfet$78_14 m1_19839_21786# vss m1_19969_21590# vss nfet$78
Xnfet$94_13 m1_13514_15478# m1_13514_15478# m1_n1927_20274# m1_n1927_20274# m1_16890_20470#
+ vss nfet$94
Xpfet$66_79 w_n11156_26804# m1_15564_15778# m1_14743_16202# m1_14482_17343# pfet$66
Xpfet$66_68 w_n11156_26804# w_n11156_26804# m1_22034_17714# m1_22493_16080# pfet$66
Xpfet$66_13 w_n11156_26804# w_n11156_26804# m1_5148_15478# sd6 pfet$66
Xpfet$66_24 w_n11156_26804# m1_6377_16202# m1_5892_17518# m1_6275_17836# pfet$66
Xpfet$66_35 w_n11156_26804# w_n11156_26804# m1_9015_17714# m1_9485_17714# pfet$66
Xpfet$66_46 w_n11156_26804# w_n11156_26804# m1_n2250_17343# m1_649_17714# pfet$66
Xpfet$66_57 w_n11156_26804# m1_n1989_16202# m1_n2474_17518# m1_n2091_17836# pfet$66
Xpfet$72_1 w_n11156_26804# w_n11156_26804# m1_21880_15478# sd2 pfet$72
Xpfet$77_12 w_n11156_26804# m1_31535_22102# w_n11156_26804# m1_3871_22513# pfet$77
Xnfet$75_15 m1_26873_21786# m1_26873_21786# m1_28490_22513# m1_28490_22513# m1_28094_21586#
+ vss nfet$75
Xnfet_22 m1_29607_24346# m1_29607_24346# vss vss m1_29089_24542# vss nfet
Xnfet_11 m1_16442_24224# m1_16442_24224# m1_16086_24542# m1_16086_24542# m1_16540_24542#
+ vss nfet
Xnfet$86_14 m1_15188_21786# m1_15188_21786# vss vss m1_14026_21586# vss nfet$86
Xpfet$66_104 w_n11156_26804# w_n11156_26804# m1_14127_16080# m1_n7513_20152# pfet$66
Xnfet$77_9 sd5 vss m1_9331_15478# vss nfet$77
Xpfet$90_12 w_n11156_26804# w_n11156_26804# m1_n6973_21481# m1_n6839_21786# pfet$90
Xnfet$89_0 m1_30256_22102# vss m1_32818_21586# vss nfet$89
Xnfet$96_1 m1_n6433_17343# m1_n4377_15778# m1_n4994_16080# vss nfet$96
Xpfet$69_13 w_n11156_26804# w_n11156_26804# m1_15188_21786# m1_14556_21786# pfet$69
Xnfet$82_7 m1_25107_21786# vss m1_32193_25858# vss nfet$82
Xnfet$75_6 m1_2384_21590# m1_2384_21590# m1_3871_22513# m1_3871_22513# m1_2843_21586#
+ vss nfet$75
Xpfet$95_0 w_n11156_26804# w_n11156_26804# m1_n5227_20152# m1_n2543_20130# pfet$95
Xnfet$101_9 m1_n3184_24224# vss m1_n3541_23922# vss nfet$101
Xpfet$69_7 w_n11156_26804# w_n11156_26804# m1_4637_21786# m1_4005_21786# pfet$69
Xpfet_105 w_n11156_26804# w_n11156_26804# m1_30888_24542# m1_28492_25858# pfet
Xpfet$74_5 w_n11156_26804# m1_32675_25947# w_n11156_26804# m1_34278_25658# pfet$74
Xpfet_69 w_n11156_26804# w_n11156_26804# m1_12875_24346# m1_n7513_20152# pfet
Xpfet_58 w_n11156_26804# w_n11156_26804# m1_23964_25662# m1_23827_25858# pfet
Xpfet_47 w_n11156_26804# w_n11156_26804# m1_15943_25858# m1_17058_24346# pfet
Xpfet$71_14 w_n11156_26804# w_n11156_26804# m1_23486_19550# m1_21564_17714# pfet$71
Xpfet_36 w_n11156_26804# w_n11156_26804# m1_8692_24346# m1_n7513_20152# pfet
Xpfet_25 w_n11156_26804# w_n11156_26804# m1_4005_21786# m1_3394_25858# pfet
Xpfet_14 w_n11156_26804# w_n11156_26804# m1_11902_25662# m1_11760_25858# pfet
Xpfet$67_4 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_9877_22102# m1_9418_21590#
+ m1_9418_21590# pfet$67
Xnfet$78_15 m1_28624_21786# vss m1_29256_21786# vss nfet$78
Xnfet$94_14 m1_22205_20152# m1_22205_20152# m1_n2543_20130# m1_n2543_20130# m1_21039_20470#
+ vss nfet$94
Xpfet$66_69 w_n11156_26804# w_n11156_26804# m1_20721_15778# m1_17851_17714# pfet$66
Xpfet$66_14 w_n11156_26804# w_n11156_26804# m1_2092_17836# m1_1933_17343# pfet$66
Xpfet$66_25 w_n11156_26804# w_n11156_26804# m1_1709_17518# m1_1119_17714# pfet$66
Xpfet$66_36 w_n11156_26804# w_n11156_26804# m1_6116_17343# m1_9015_17714# pfet$66
Xpfet$66_47 w_n11156_26804# m1_11738_16080# m1_11271_18030# m1_10299_17343# pfet$66
Xpfet$66_58 w_n11156_26804# w_n11156_26804# m1_n3534_17714# m1_n3064_17714# pfet$66
Xpfet$72_2 w_n11156_26804# w_n11156_26804# m1_26063_15478# sd1 pfet$72
Xpfet$77_13 w_n11156_26804# w_n11156_26804# m1_31535_22102# m1_354_22513# pfet$77
Xnfet$75_16 m1_27003_21590# m1_27003_21590# m1_28490_22513# m1_28490_22513# m1_27462_21586#
+ vss nfet$75
Xnfet_23 m1_25424_24346# m1_25424_24346# m1_24309_25858# m1_24309_25858# m1_26371_25502#
+ vss nfet
Xnfet_12 m1_17058_24346# m1_17058_24346# m1_15943_25858# m1_15943_25858# m1_18005_25502#
+ vss nfet
Xnfet$86_15 m1_14556_21786# m1_14556_21786# vss vss m1_13394_21586# vss nfet$86
Xpfet$66_105 w_n11156_26804# w_n11156_26804# m1_14258_17518# m1_13668_17714# pfet$66
Xpfet$90_13 w_n11156_26804# w_n11156_26804# m1_n6839_21786# m1_n6380_21786# pfet$90
Xnfet$89_1 m1_31535_22102# m1_32818_21586# vss vss nfet$89
Xnfet$96_2 m1_n6274_17836# m1_n5351_15778# m1_n6172_16202# vss nfet$96
Xnfet$82_8 m1_32193_25858# vss m1_32330_25662# vss nfet$82
Xpfet$69_14 w_n11156_26804# w_n11156_26804# m1_19969_21590# m1_19839_21786# pfet$69
Xnfet$75_7 m1_5771_21786# m1_5771_21786# m1_7388_22513# m1_7388_22513# m1_6992_21586#
+ vss nfet$75
Xpfet$69_8 w_n11156_26804# w_n11156_26804# m1_2384_21590# m1_2254_21786# pfet$69
Xpfet$95_1 w_n11156_26804# m1_n4485_20152# w_n11156_26804# m1_n3206_20274# pfet$95
Xpfet$88_0 w_n11156_26804# w_n11156_26804# m1_n7320_25516# m1_n7186_25858# pfet$88
Xpfet$74_6 w_n11156_26804# w_n11156_26804# m1_32818_24542# m1_33174_24224# pfet$74
Xpfet_59 w_n11156_26804# w_n11156_26804# m1_16322_21786# pd6 pfet
Xpfet_48 w_n11156_26804# m1_16085_25662# m1_15822_23922# m1_15598_25662# pfet
Xpfet$71_15 w_n11156_26804# w_n11156_26804# m1_22205_20152# m1_17697_15478# pfet$71
Xpfet_37 w_n11156_26804# w_n11156_26804# m1_9973_24542# m1_7577_25858# pfet
Xpfet_26 w_n11156_26804# m1_4997_25658# m1_5790_24542# m1_3049_25662# pfet
Xpfet_15 w_n11156_26804# m1_11902_25662# m1_11639_23922# m1_11415_25662# pfet
Xnfet$106_0 m1_n6839_20152# vss m1_n8145_21908# vss nfet$106
Xpfet_106 w_n11156_26804# w_n11156_26804# m1_25107_21786# m1_28492_25858# pfet
Xnfet$78_16 m1_26873_21786# vss m1_27003_21590# vss nfet$78
Xpfet$67_5 w_n11156_26804# m1_9645_21447# m1_9645_21447# m1_9877_22102# m1_11671_21786#
+ m1_11671_21786# pfet$67
Xnfet$94_15 m1_17697_15478# m1_17697_15478# m1_n2543_20130# m1_n2543_20130# m1_20407_20470#
+ vss nfet$94
Xpfet$66_15 w_n11156_26804# w_n11156_26804# m1_5302_17714# m1_5761_16080# pfet$66
Xpfet$66_26 w_n11156_26804# w_n11156_26804# m1_4832_17714# m1_5302_17714# pfet$66
Xpfet$66_37 w_n11156_26804# m1_7555_16080# m1_7088_18030# m1_6116_17343# pfet$66
Xpfet$66_48 w_n11156_26804# w_n11156_26804# m1_n3064_17714# m1_n2605_16080# pfet$66
Xpfet$66_59 w_n11156_26804# w_n11156_26804# m1_n2605_16080# m1_n7513_20152# pfet$66
Xnfet$75_17 m1_12935_21590# m1_12935_21590# m1_14422_22513# m1_14422_22513# m1_13394_21586#
+ vss nfet$75
Xpfet$70_0 w_n11156_26804# w_n11156_26804# m1_n6274_17836# m1_n6433_17343# pfet$70
Xnfet_24 m1_30095_25658# m1_30095_25658# vss vss m1_30554_25502# vss nfet
Xnfet_13 m1_13363_25658# m1_13363_25658# vss vss m1_13822_25502# vss nfet
Xpfet$66_106 w_n11156_26804# w_n11156_26804# m1_14482_17343# m1_17381_17714# pfet$66
Xnfet$86_16 m1_28624_21786# m1_28624_21786# vss vss m1_27462_21586# vss nfet$86
Xnfet$96_3 m1_n6433_17343# m1_n6172_16202# m1_n6657_17518# vss nfet$96
Xnfet$82_9 m1_n7513_20152# vss m1_33790_24346# vss nfet$82
Xpfet$69_15 w_n11156_26804# w_n11156_26804# m1_27003_21590# m1_26873_21786# pfet$69
Xpfet$69_9 w_n11156_26804# w_n11156_26804# m1_22222_21786# m1_21590_21786# pfet$69
Xnfet$75_8 m1_23486_21590# m1_23486_21590# m1_24973_22513# m1_24973_22513# m1_23945_21586#
+ vss nfet$75
Xnfet$94_0 m1_4620_20152# m1_4620_20152# m1_2590_19404# m1_2590_19404# m1_3454_20470#
+ vss nfet$94
Xpfet$95_2 w_n11156_26804# m1_n6839_20152# w_n11156_26804# m1_n927_19404# pfet$95
Xpfet$88_1 w_n11156_26804# w_n11156_26804# m1_n6111_25858# m1_n6856_24542# pfet$88
Xpfet$71_16 w_n11156_26804# w_n11156_26804# m1_19969_19550# m1_17381_17714# pfet$71
Xnfet$106_1 m1_n5227_20152# vss m1_n6380_21786# vss nfet$106
Xpfet_107 w_n11156_26804# m1_24309_25858# w_n11156_26804# m1_25912_25658# pfet
Xpfet$74_7 w_n11156_26804# m1_32818_24542# w_n11156_26804# m1_33790_24346# pfet$74
Xpfet_49 w_n11156_26804# m1_20126_25858# w_n11156_26804# m1_21729_25658# pfet
Xpfet_38 w_n11156_26804# w_n11156_26804# m1_16085_25662# m1_15943_25858# pfet
Xpfet_27 w_n11156_26804# w_n11156_26804# m1_11278_25858# m1_7522_21786# pfet
Xpfet_16 w_n11156_26804# w_n11156_26804# m1_5771_21786# pd3 pfet
Xpfet$67_6 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_10505_22402# m1_9288_21786#
+ m1_9288_21786# pfet$67
Xnfet$78_17 m1_25107_21786# vss m1_25739_21786# vss nfet$78
Xnfet$94_16 m1_25722_20152# m1_25722_20152# m1_n3206_20274# m1_n3206_20274# m1_24556_20470#
+ vss nfet$94
Xpfet$66_16 w_n11156_26804# w_n11156_26804# m1_3989_15778# m1_1119_17714# pfet$66
Xpfet$66_27 w_n11156_26804# m1_2194_16202# m1_1709_17518# m1_2092_17836# pfet$66
Xpfet$66_38 w_n11156_26804# w_n11156_26804# m1_7088_18030# m1_7198_15778# pfet$66
Xpfet$66_49 w_n11156_26804# m1_n194_15778# m1_n811_16080# m1_n2091_17836# pfet$66
Xpfet$70_1 w_n11156_26804# w_n11156_26804# m1_n4377_15778# m1_n7247_17714# pfet$70
Xnfet$101_10 vss vss m1_n4978_24224# vss nfet$101
Xpfet$66_107 w_n11156_26804# m1_15921_16080# m1_15454_18030# m1_14482_17343# pfet$66
Xnfet_25 m1_29607_24346# m1_29607_24346# m1_28492_25858# m1_28492_25858# m1_30554_25502#
+ vss nfet
Xnfet$86_17 m1_29256_21786# m1_29256_21786# vss vss m1_28094_21586# vss nfet$86
Xnfet_14 m1_12875_24346# m1_12875_24346# m1_11760_25858# m1_11760_25858# m1_13822_25502#
+ vss nfet
Xnfet$96_4 m1_27031_17343# m1_27292_16202# m1_26807_17518# vss nfet$96
Xpfet$69_16 w_n11156_26804# w_n11156_26804# m1_29256_21786# m1_28624_21786# pfet$69
Xnfet$75_9 m1_23356_21786# m1_23356_21786# m1_24973_22513# m1_24973_22513# m1_24577_21586#
+ vss nfet$75
Xnfet$87_0 m1_21456_22513# m1_21456_22513# m1_30256_19792# m1_30256_19792# m1_30492_20470#
+ vss nfet$87
Xnfet$94_1 m1_1103_20152# m1_1103_20152# m1_n927_19404# m1_n927_19404# m1_n63_20470#
+ vss nfet$94
Xpfet$95_3 w_n11156_26804# m1_n5227_20152# w_n11156_26804# m1_n1927_20274# pfet$95
Xpfet$71_17 w_n11156_26804# w_n11156_26804# m1_25722_20152# m1_21880_15478# pfet$71
Xnfet$106_2 m1_n4485_20152# m1_n6380_21786# vss vss nfet$106
Xpfet_108 w_n11156_26804# w_n11156_26804# m1_25424_24346# m1_n7513_20152# pfet
Xpfet_39 w_n11156_26804# w_n11156_26804# m1_15598_25662# m1_15461_25858# pfet
Xpfet_28 w_n11156_26804# m1_11639_23922# m1_11903_24542# m1_11278_25858# pfet
Xpfet_17 w_n11156_26804# w_n11156_26804# m1_7577_25858# m1_8692_24346# pfet
Xpfet$67_7 w_n11156_26804# m1_354_22513# m1_354_22513# m1_n674_22102# m1_1120_21786#
+ m1_1120_21786# pfet$67
Xnfet$94_17 m1_21880_15478# m1_21880_15478# m1_n3206_20274# m1_n3206_20274# m1_23924_20470#
+ vss nfet$94
Xpfet$93_0 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_n8047_19550# m1_n7513_20152#
+ m1_n7513_20152# pfet$93
Xpfet$66_17 w_n11156_26804# w_n11156_26804# m1_n2091_17836# m1_n2250_17343# pfet$66
Xpfet$66_28 w_n11156_26804# m1_2905_18030# w_n11156_26804# m1_1578_16080# pfet$66
Xpfet$66_39 w_n11156_26804# m1_7088_18030# w_n11156_26804# m1_5761_16080# pfet$66
Xpfet$70_2 w_n11156_26804# w_n11156_26804# m1_n5351_15778# m1_n4994_16080# pfet$70
Xnfet$101_11 m1_n10452_25858# vss m1_n4847_25662# vss nfet$101
Xnfet_26 m1_25912_25658# m1_25912_25658# vss vss m1_26371_25502# vss nfet
Xnfet_15 m1_25424_24346# m1_25424_24346# vss vss m1_24906_24542# vss nfet
Xpfet$66_108 w_n11156_26804# w_n11156_26804# m1_15454_18030# m1_15564_15778# pfet$66
Xnfet$96_5 m1_27031_17343# m1_29087_15778# m1_28470_16080# vss nfet$96
Xpfet$69_17 w_n11156_26804# w_n11156_26804# m1_25739_21786# m1_25107_21786# pfet$69
Xnfet$87_1 m1_24973_22513# m1_24973_22513# vss vss m1_30492_20470# vss nfet$87
Xnfet$94_2 m1_n3218_15478# m1_n3218_15478# m1_2590_19404# m1_2590_19404# m1_2822_20470#
+ vss nfet$94
Xpfet$95_4 w_n11156_26804# w_n11156_26804# m1_n4485_20152# m1_n3822_20130# pfet$95
Xnfet$106_3 m1_n5227_21418# vss m1_n5764_21786# vss nfet$106
Xpfet_109 w_n11156_26804# m1_12259_24224# m1_13363_25658# m1_11278_25858# pfet
Xpfet_29 w_n11156_26804# w_n11156_26804# m1_11903_24542# m1_12259_24224# pfet
Xpfet_18 w_n11156_26804# w_n11156_26804# m1_11415_25662# m1_11278_25858# pfet
Xpfet$67_8 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_6360_22102# m1_5901_21590#
+ m1_5901_21590# pfet$67
Xpfet$93_1 w_n11156_26804# m1_n8283_19850# m1_n8283_19850# m1_n8047_19550# m1_n8283_20611#
+ m1_n8283_20611# pfet$93
Xpfet$86_0 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_n6624_23622# m1_n7082_23622#
+ m1_n7082_23622# pfet$86
Xpfet$66_18 w_n11156_26804# m1_1119_17714# w_n11156_26804# m1_2194_16202# pfet$66
Xpfet$66_29 w_n11156_26804# w_n11156_26804# m1_1578_16080# m1_n7513_20152# pfet$66
Xnfet$104_0 m1_n7186_25858# vss m1_n7320_25516# vss nfet$104
Xpfet$70_3 w_n11156_26804# w_n11156_26804# m1_n6657_17518# m1_n7247_17714# pfet$70
Xnfet$101_12 m1_n10452_25858# vss m1_n5571_25662# vss nfet$101
Xnfet_27 m1_12875_24346# m1_12875_24346# vss vss m1_12357_24542# vss nfet
Xpfet$66_109 w_n11156_26804# w_n11156_26804# m1_10299_17343# m1_13198_17714# pfet$66
Xnfet_16 m1_24808_24224# m1_24808_24224# m1_24452_24542# m1_24452_24542# m1_24906_24542#
+ vss nfet
Xnfet$96_6 m1_27190_17836# m1_28113_15778# m1_27292_16202# vss nfet$96
Xpfet$95_5 w_n11156_26804# w_n11156_26804# m1_n6839_20152# m1_n6973_21481# pfet$95
Xnfet$87_2 m1_14422_22513# m1_14422_22513# m1_31535_19792# m1_31535_19792# m1_31771_20470#
+ vss nfet$87
Xnfet$94_3 m1_8137_20152# m1_8137_20152# m1_6107_19404# m1_6107_19404# m1_6971_20470#
+ vss nfet$94
Xnfet$106_4 m1_n4485_21904# m1_n5764_21786# vss vss nfet$106
Xpfet_19 w_n11156_26804# w_n11156_26804# m1_7095_25858# m1_4005_21786# pfet
Xpfet$67_9 w_n11156_26804# m1_3871_22513# m1_3871_22513# m1_3471_22402# m1_4005_21786#
+ m1_4005_21786# pfet$67
Xnfet$92_0 fout vss m1_35837_22102# vss nfet$92
Xpfet$93_2 w_n11156_26804# m1_n8283_20611# m1_n8283_20611# m1_n8047_22344# m1_n8145_21908#
+ m1_n8145_21908# pfet$93
Xpfet$79_0 w_n11156_26804# m1_n647_25662# m1_n910_23922# m1_n1134_25662# pfet$79
Xpfet$86_1 w_n11156_26804# m1_n6856_24542# m1_n6856_24542# m1_n6624_23622# m1_n8283_19850#
+ m1_n8283_19850# pfet$86
Xpfet$66_19 w_n11156_26804# m1_3015_15778# m1_2194_16202# m1_1933_17343# pfet$66
Xnfet$104_1 m1_n6856_24542# vss m1_n6111_25858# vss nfet$104
Xpfet$70_4 w_n11156_26804# w_n11156_26804# m1_n6433_17343# m1_n3534_17714# pfet$70
Xnfet$101_13 fin vss m1_n4623_25487# vss nfet$101
Xnfet_17 m1_20625_24224# m1_20625_24224# m1_20269_24542# m1_20269_24542# m1_20723_24542#
+ vss nfet
Xnfet$96_7 m1_27190_17836# m1_28470_16080# m1_28003_18030# vss nfet$96
Xnfet$87_3 m1_17939_22513# m1_17939_22513# vss vss m1_31771_20470# vss nfet$87
Xnfet$94_4 m1_965_15478# m1_965_15478# m1_6107_19404# m1_6107_19404# m1_6339_20470#
+ vss nfet$94
Xnfet$106_5 m1_n6839_21786# vss m1_n6973_21481# vss nfet$106
Xnfet$92_1 define m1_35837_22102# vss vss nfet$92
Xpfet$93_3 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_n8047_22344# m1_n8283_19850#
+ m1_n8283_19850# pfet$93
Xnfet$85_0 m1_n290_24224# m1_n290_24224# m1_n646_24542# m1_n646_24542# m1_n192_24542#
+ vss nfet$85
Xpfet$79_1 w_n11156_26804# m1_n910_23922# m1_n646_24542# m1_n1271_25858# pfet$79
Xpfet$91_0 w_n11156_26804# w_n11156_26804# m1_n10796_25662# m1_n10933_25858# pfet$91
Xpfet$67_30 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_17539_22402# m1_16322_21786#
+ m1_16322_21786# pfet$67
Xpfet$70_5 w_n11156_26804# w_n11156_26804# m1_n6788_16080# m1_n7513_20152# pfet$70
Xnfet$81_10 m1_26217_17714# vss m1_29087_15778# vss nfet$81
Xnfet_18 m1_21241_24346# m1_21241_24346# vss vss m1_20723_24542# vss nfet
Xnfet$76_10 m1_9015_17714# m1_9015_17714# vss vss m1_14005_20470# vss nfet$76
Xnfet$87_4 m1_32818_20470# m1_32818_20470# vss vss m1_34329_20470# vss nfet$87
Xnfet$94_5 m1_5148_15478# m1_5148_15478# m1_9624_19404# m1_9624_19404# m1_9856_20470#
+ vss nfet$94
Xnfet$85_1 m1_814_25658# m1_814_25658# vss vss m1_1273_25502# vss nfet$85
Xpfet$79_2 w_n11156_26804# m1_n290_24224# m1_814_25658# m1_n1271_25858# pfet$79
Xnfet$78_0 m1_n1263_21786# vss m1_n1133_21590# vss nfet$78
Xpfet$84_0 w_n11156_26804# m1_n4377_15778# m1_n4994_16080# m1_n6274_17836# pfet$84
Xpfet$91_1 w_n11156_26804# w_n11156_26804# m1_n10309_25662# m1_n10452_25858# pfet$91
Xnfet$79_10 m1_26063_15478# vss m1_29239_20152# vss nfet$79
Xnfet$102_0 m1_n9952_24224# m1_n9952_24224# m1_n10308_24542# m1_n10308_24542# m1_n9854_24542#
+ vss nfet$102
Xpfet$67_31 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_27462_22102# m1_27003_21590#
+ m1_27003_21590# pfet$67
Xpfet$67_20 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_20428_22102# m1_19969_21590#
+ m1_19969_21590# pfet$67
Xpfet$70_6 w_n11156_26804# w_n11156_26804# m1_n7383_17599# m1_n7247_17714# pfet$70
Xnfet$81_11 m1_27031_17343# vss m1_27190_17836# vss nfet$81
Xnfet_19 m1_21729_25658# m1_21729_25658# vss vss m1_22188_25502# vss nfet
Xnfet$76_11 m1_13198_17714# m1_13198_17714# vss vss m1_17522_20470# vss nfet$76
Xnfet$87_10 m1_354_22513# m1_354_22513# m1_31535_22102# m1_31535_22102# m1_31771_21430#
+ vss nfet$87
Xnfet$87_5 m1_32818_21586# m1_32818_21586# m1_34093_19792# m1_34093_19792# m1_34329_20470#
+ vss nfet$87
Xnfet$94_6 m1_11654_20152# m1_11654_20152# m1_9624_19404# m1_9624_19404# m1_10488_20470#
+ vss nfet$94
Xpfet$79_3 w_n11156_26804# m1_814_25658# m1_1607_24542# m1_n1134_25662# pfet$79
Xnfet$85_2 m1_326_24346# m1_326_24346# m1_n789_25858# m1_n789_25858# m1_1273_25502#
+ vss nfet$85
Xnfet$78_1 m1_11039_21786# vss m1_11671_21786# vss nfet$78
Xnfet$90_0 m1_34093_19792# vss m1_34843_21786# vss nfet$90
Xpfet$77_0 w_n11156_26804# m1_31535_19792# w_n11156_26804# m1_17939_22513# pfet$77
Xpfet$84_1 w_n11156_26804# m1_n5351_15778# m1_n6172_16202# m1_n6433_17343# pfet$84
Xpfet$91_2 w_n11156_26804# w_n11156_26804# m1_n9952_24224# m1_n10572_23922# pfet$91
Xnfet$79_11 m1_9331_15478# vss m1_15171_20152# vss nfet$79
Xnfet$102_1 m1_n9336_24346# m1_n9336_24346# m1_n8625_26174# m1_n8625_26174# m1_n8389_25502#
+ vss nfet$102
Xpfet$67_32 w_n11156_26804# m1_28490_22513# m1_28490_22513# m1_28090_22402# m1_28624_21786#
+ m1_28624_21786# pfet$67
Xpfet$67_21 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_21056_22402# m1_19839_21786#
+ m1_19839_21786# pfet$67
Xpfet$70_7 w_n11156_26804# w_n11156_26804# m1_27190_17836# m1_27031_17343# pfet$70
Xpfet$67_10 w_n11156_26804# m1_3871_22513# m1_3871_22513# m1_2843_22102# m1_4637_21786#
+ m1_4637_21786# pfet$67
Xnfet$81_12 m1_28470_16080# vss m1_28113_15778# vss nfet$81
Xnfet$76_12 m1_16452_19550# m1_16452_19550# vss vss m1_16890_20470# vss nfet$76
Xnfet$87_11 m1_3871_22513# m1_3871_22513# vss vss m1_31771_21430# vss nfet$87
Xnfet$87_6 m1_28490_22513# m1_28490_22513# vss vss m1_34329_21430# vss nfet$87
Xnfet$94_7 m1_n7401_15478# m1_n7401_15478# m1_n927_19404# m1_n927_19404# m1_n695_20470#
+ vss nfet$94
Xpfet$79_4 w_n11156_26804# m1_33174_24224# m1_34278_25658# m1_32193_25858# pfet$79
Xnfet$85_3 m1_326_24346# m1_326_24346# vss vss m1_n192_24542# vss nfet$85
Xnfet$78_2 m1_12805_21786# vss m1_12935_21590# vss nfet$78
Xpfet$91_3 w_n11156_26804# w_n11156_26804# m1_n4978_24224# vss pfet$91
Xnfet$79_12 m1_13514_15478# vss m1_18688_20152# vss nfet$79
Xnfet$90_1 m1_30256_19792# vss m1_32818_20470# vss nfet$90
Xpfet$77_1 w_n11156_26804# w_n11156_26804# m1_30256_19792# m1_21456_22513# pfet$77
Xpfet$84_2 w_n11156_26804# m1_n4994_16080# m1_n5461_18030# m1_n6433_17343# pfet$84
Xnfet$102_2 m1_n8848_25658# m1_n8848_25658# vss vss m1_n8389_25502# vss nfet$102
Xnfet$83_0 m1_n1134_25662# m1_n910_23922# m1_n646_24542# vss nfet$83
Xpfet$67_33 w_n11156_26804# m1_28490_22513# m1_28490_22513# m1_27462_22102# m1_29256_21786#
+ m1_29256_21786# pfet$67
Xpfet$67_22 w_n11156_26804# m1_21456_22513# m1_21456_22513# m1_20428_22102# m1_22222_21786#
+ m1_22222_21786# pfet$67
Xpfet$70_8 w_n11156_26804# w_n11156_26804# m1_28113_15778# m1_28470_16080# pfet$70
Xpfet$67_11 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_2843_22102# m1_2384_21590#
+ m1_2384_21590# pfet$67
Xnfet$81_13 m1_26217_17714# vss m1_25747_17714# vss nfet$81
Xnfet$76_13 m1_19969_19550# m1_19969_19550# vss vss m1_20407_20470# vss nfet$76
Xnfet$87_7 m1_34843_21786# m1_34843_21786# m1_34093_22102# m1_34093_22102# m1_34329_21430#
+ vss nfet$87
Xnfet$94_8 m1_26063_15478# m1_26063_15478# m1_n3822_20130# m1_n3822_20130# m1_27441_20470#
+ vss nfet$94
Xpfet$91_10 w_n11156_26804# w_n11156_26804# m1_n10933_25858# fin pfet$91
Xpfet$79_5 w_n11156_26804# m1_32817_25662# m1_32554_23922# m1_32330_25662# pfet$79
Xnfet$85_4 m1_33174_24224# m1_33174_24224# m1_32818_24542# m1_32818_24542# m1_33272_24542#
+ vss nfet$85
Xnfet$78_3 m1_9288_21786# vss m1_9418_21590# vss nfet$78
Xnfet$90_2 m1_31535_19792# m1_32818_20470# vss vss nfet$90
Xpfet$77_2 w_n11156_26804# m1_30256_19792# w_n11156_26804# m1_24973_22513# pfet$77
Xnfet$76_0 m1_n3534_17714# m1_n3534_17714# vss vss m1_3454_20470# vss nfet$76
Xpfet$84_3 w_n11156_26804# m1_n6172_16202# m1_n6657_17518# m1_n6274_17836# pfet$84
Xpfet$91_4 w_n11156_26804# w_n11156_26804# m1_n5571_25662# m1_n10452_25858# pfet$91
Xnfet$83_1 m1_n1271_25858# m1_n647_25662# m1_n910_23922# vss nfet$83
Xpfet$67_34 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_28090_22402# m1_26873_21786#
+ m1_26873_21786# pfet$67
Xpfet$67_23 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_23945_22102# m1_23486_21590#
+ m1_23486_21590# pfet$67
Xnfet$79_13 m1_13198_17714# vss m1_16452_19550# vss nfet$79
Xpfet$67_12 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_3471_22402# m1_2254_21786#
+ m1_2254_21786# pfet$67
Xnfet$102_3 m1_n9336_24346# m1_n9336_24346# vss vss m1_n9854_24542# vss nfet$102
Xpfet$82_0 w_n11156_26804# w_n11156_26804# fout m1_34093_22102# pfet$82
Xpfet$70_9 w_n11156_26804# w_n11156_26804# m1_29087_15778# m1_26217_17714# pfet$70
Xnfet$100_0 m1_n927_19404# m1_n927_19404# vss vss m1_n6282_20470# vss nfet$100
Xnfet$76_14 m1_17381_17714# m1_17381_17714# vss vss m1_21039_20470# vss nfet$76
Xnfet$87_8 m1_9645_21447# m1_9645_21447# vss vss m1_30492_21430# vss nfet$87
Xnfet$94_9 m1_29239_20152# m1_29239_20152# m1_n3822_20130# m1_n3822_20130# m1_28073_20470#
+ vss nfet$94
Xpfet$91_11 w_n11156_26804# w_n11156_26804# m1_n9336_24346# vss pfet$91
Xnfet_0 m1_4509_24346# m1_4509_24346# vss vss m1_3991_24542# vss nfet
Xpfet$79_6 w_n11156_26804# m1_34278_25658# m1_35071_24542# m1_32330_25662# pfet$79
Xnfet$85_5 m1_33790_24346# m1_33790_24346# vss vss m1_33272_24542# vss nfet$85
Xnfet$78_4 m1_7522_21786# vss m1_8154_21786# vss nfet$78
Xnfet$74_80 m1_28147_25662# m1_28991_24224# m1_30095_25658# vss nfet$74
Xnfet$90_3 m1_34093_22102# vss fout vss nfet$90
Xpfet$77_3 w_n11156_26804# w_n11156_26804# m1_34843_21786# m1_34093_19792# pfet$77
Xpfet$84_4 w_n11156_26804# m1_28113_15778# m1_27292_16202# m1_27031_17343# pfet$84
Xnfet$83_2 m1_n1271_25858# m1_814_25658# m1_1607_24542# vss nfet$83
Xnfet$76_1 m1_2384_19550# m1_2384_19550# vss vss m1_2822_20470# vss nfet$76
Xpfet$91_5 w_n11156_26804# w_n11156_26804# m1_n4847_25662# m1_n10452_25858# pfet$91
Xnfet$79_14 m1_21564_17714# vss m1_23486_19550# vss nfet$79
Xnfet$102_4 m1_n4978_24224# m1_n4978_24224# m1_n10452_25858# m1_n10452_25858# m1_n4880_24542#
+ vss nfet$102
Xpfet$67_35 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_13394_22102# m1_12935_21590#
+ m1_12935_21590# pfet$67
Xpfet$67_24 w_n11156_26804# m1_17939_22513# m1_17939_22513# m1_16911_22102# m1_18705_21786#
+ m1_18705_21786# pfet$67
Xpfet$67_13 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_6988_22402# m1_5771_21786#
+ m1_5771_21786# pfet$67
Xpfet$75_0 w_n11156_26804# m1_32818_21586# m1_32818_21586# m1_33050_22344# m1_30256_22102#
+ m1_30256_22102# pfet$75
Xnfet$100_1 m1_n3822_20130# m1_n3822_20130# m1_n4485_20152# m1_n4485_20152# m1_n3724_20470#
+ vss nfet$100
Xnfet$76_15 m1_21564_17714# m1_21564_17714# vss vss m1_24556_20470# vss nfet$76
Xnfet$87_9 m1_7388_22513# m1_7388_22513# m1_30256_22102# m1_30256_22102# m1_30492_21430#
+ vss nfet$87
Xnfet$77_80 m1_18824_17836# m1_19747_15778# m1_18926_16202# vss nfet$77
Xpfet$91_12 w_n11156_26804# w_n11156_26804# m1_n7082_23622# m1_n8625_26174# pfet$91
Xnfet$99_0 m1_n7082_23622# m1_n6856_24542# vss vss nfet$99
Xnfet_1 m1_3893_24224# m1_3893_24224# m1_3537_24542# m1_3537_24542# m1_3991_24542#
+ vss nfet
Xpfet$79_7 w_n11156_26804# m1_32554_23922# m1_32818_24542# m1_32193_25858# pfet$79
Xnfet$85_6 m1_33790_24346# m1_33790_24346# m1_32675_25947# m1_32675_25947# m1_34737_25502#
+ vss nfet$85
Xnfet$78_5 m1_488_21786# vss m1_1120_21786# vss nfet$78
Xnfet$74_81 m1_n7513_20152# vss m1_25424_24346# vss nfet$74
Xnfet$74_70 m1_21590_21786# vss m1_28010_25858# vss nfet$74
Xnfet$90_4 m1_31535_22102# m1_32818_21586# vss vss nfet$90
Xpfet$77_4 w_n11156_26804# m1_34093_19792# w_n11156_26804# m1_32818_20470# pfet$77
Xpfet$84_5 w_n11156_26804# m1_29087_15778# m1_28470_16080# m1_27190_17836# pfet$84
Xnfet$83_3 m1_n1134_25662# m1_n290_24224# m1_814_25658# vss nfet$83
Xnfet$76_2 m1_5901_19550# m1_5901_19550# vss vss m1_6339_20470# vss nfet$76
Xpfet$91_6 w_n11156_26804# w_n11156_26804# m1_n4623_25487# fin pfet$91
Xnfet$79_15 m1_17697_15478# vss m1_22205_20152# vss nfet$79
Xnfet$102_5 m1_n4362_24346# m1_n4362_24346# vss vss m1_n4880_24542# vss nfet$102
Xpfet$67_25 w_n11156_26804# m1_17939_22513# m1_17939_22513# m1_17539_22402# m1_18073_21786#
+ m1_18073_21786# pfet$67
Xpfet$67_14 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_n46_22402# m1_n1263_21786#
+ m1_n1263_21786# pfet$67
Xpfet$75_1 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_33050_22344# m1_31535_22102#
+ m1_31535_22102# pfet$75
Xpfet$68_0 w_n11156_26804# m1_2590_19404# m1_2590_19404# m1_3458_19550# m1_n3534_17714#
+ m1_n3534_17714# pfet$68
Xnfet$81_0 m1_n3534_17714# vss m1_n6433_17343# vss nfet$81
Xnfet$100_2 m1_n2543_20130# m1_n2543_20130# m1_n5227_20152# m1_n5227_20152# m1_n2445_20470#
+ vss nfet$100
Xnfet$76_16 m1_23486_19550# m1_23486_19550# vss vss m1_23924_20470# vss nfet$76
Xnfet$77_81 m1_13198_17714# vss m1_10299_17343# vss nfet$77
Xnfet$77_70 m1_n7513_20152# vss m1_18310_16080# vss nfet$77
Xpfet$91_13 w_n11156_26804# w_n11156_26804# m1_n8055_24542# m1_n8625_26174# pfet$91
Xnfet$99_1 m1_n8283_19850# vss m1_n6856_24542# vss nfet$99
Xnfet_2 m1_4997_25658# m1_4997_25658# vss vss m1_5456_25502# vss nfet
Xnfet$85_7 m1_34278_25658# m1_34278_25658# vss vss m1_34737_25502# vss nfet$85
Xnfet$78_6 m1_5771_21786# vss m1_5901_21590# vss nfet$78
Xnfet$74_82 m1_11415_25662# m1_12259_24224# m1_13363_25658# vss nfet$74
Xnfet$74_71 m1_28147_25662# m1_28371_23922# m1_28635_24542# vss nfet$74
Xnfet$90_5 m1_30256_22102# vss m1_32818_21586# vss nfet$90
Xnfet$74_60 pd6 vss m1_16322_21786# vss nfet$74
Xpfet$84_6 w_n11156_26804# m1_28470_16080# m1_28003_18030# m1_27031_17343# pfet$84
Xpfet$77_5 w_n11156_26804# w_n11156_26804# m1_34093_19792# m1_32818_21586# pfet$77
Xpfet$91_7 w_n11156_26804# w_n11156_26804# m1_n3541_23922# m1_n3184_24224# pfet$91
Xnfet$83_4 m1_32193_25858# m1_34278_25658# m1_35071_24542# vss nfet$83
Xnfet$79_16 m1_17381_17714# vss m1_19969_19550# vss nfet$79
Xnfet$76_3 m1_4832_17714# m1_4832_17714# vss vss m1_10488_20470# vss nfet$76
Xnfet$102_6 m1_n4978_24224# m1_n4978_24224# vss vss m1_n3415_25502# vss nfet$102
Xpfet$67_26 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_16911_22102# m1_16452_21590#
+ m1_16452_21590# pfet$67
Xpfet$67_15 w_n11156_26804# m1_354_22513# m1_354_22513# m1_n46_22402# m1_488_21786#
+ m1_488_21786# pfet$67
Xnfet$74_0 m1_3394_25858# vss m1_5790_24542# vss nfet$74
Xpfet$68_1 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_2822_19850# m1_4620_20152#
+ m1_4620_20152# pfet$68
Xnfet$81_1 m1_n7513_20152# vss m1_n6788_16080# vss nfet$81
Xnfet$100_3 m1_n1927_20274# m1_n1927_20274# vss vss m1_n2445_20470# vss nfet$100
Xnfet$76_17 m1_12935_19550# m1_12935_19550# vss vss m1_13373_20470# vss nfet$76
Xpfet$80_0 w_n11156_26804# w_n11156_26804# m1_n1263_21786# pd1 pfet$80
Xnfet$77_82 m1_10299_17343# vss m1_10458_17836# vss nfet$77
Xnfet$77_71 m1_14641_17836# m1_15921_16080# m1_15454_18030# vss nfet$77
Xnfet$77_60 m1_18665_17343# vss m1_18824_17836# vss nfet$77
Xnfet_3 m1_4509_24346# m1_4509_24346# m1_3394_25858# m1_3394_25858# m1_5456_25502#
+ vss nfet
Xnfet$78_7 m1_4005_21786# vss m1_4637_21786# vss nfet$78
Xnfet$74_72 m1_23827_25858# m1_25912_25658# m1_26705_24542# vss nfet$74
Xnfet$74_61 m1_23964_25662# m1_24808_24224# m1_25912_25658# vss nfet$74
Xnfet$74_50 m1_n7513_20152# vss m1_21241_24346# vss nfet$74
Xnfet$109_0 m1_n6839_20152# vss m1_n8145_21908# vss nfet$109
Xpfet$91_8 w_n11156_26804# w_n11156_26804# m1_n2567_23922# m1_n7320_25516# pfet$91
Xnfet$79_17 m1_21880_15478# vss m1_25722_20152# vss nfet$79
Xnfet$83_5 m1_32330_25662# m1_33174_24224# m1_34278_25658# vss nfet$83
Xpfet$84_7 w_n11156_26804# m1_27292_16202# m1_26807_17518# m1_27190_17836# pfet$84
Xpfet$77_6 w_n11156_26804# w_n11156_26804# m1_31535_19792# m1_14422_22513# pfet$77
Xnfet$76_4 m1_9418_19550# m1_9418_19550# vss vss m1_9856_20470# vss nfet$76
Xnfet$102_7 m1_n3541_23922# m1_n3541_23922# m1_n3651_26174# m1_n3651_26174# m1_n3415_25502#
+ vss nfet$102
Xpfet$67_27 w_n11156_26804# m1_14422_22513# m1_14422_22513# m1_14022_22402# m1_14556_21786#
+ m1_14556_21786# pfet$67
Xpfet$67_16 w_n11156_26804# m1_24973_22513# m1_24973_22513# m1_23945_22102# m1_25739_21786#
+ m1_25739_21786# pfet$67
Xnfet$74_1 m1_2912_25858# m1_4997_25658# m1_5790_24542# vss nfet$74
Xpfet$68_2 w_n11156_26804# m1_2590_19404# m1_2590_19404# m1_2822_19850# m1_2384_19550#
+ m1_2384_19550# pfet$68
Xnfet$81_2 m1_n4994_16080# vss m1_n5351_15778# vss nfet$81
Xnfet$100_4 m1_n3206_20274# m1_n3206_20274# vss vss m1_n3724_20470# vss nfet$100
Xpfet$80_1 w_n11156_26804# w_n11156_26804# m1_2254_21786# pd2 pfet$80
Xpfet$73_0 w_n11156_26804# w_n11156_26804# m1_n647_25662# m1_n789_25858# pfet$73
Xnfet$77_72 m1_17851_17714# vss m1_18441_17518# vss nfet$77
Xnfet$77_61 m1_20104_16080# vss m1_19747_15778# vss nfet$77
Xnfet$77_50 m1_25747_17714# vss m1_22848_17343# vss nfet$77
Xnfet_4 m1_12259_24224# m1_12259_24224# m1_11903_24542# m1_11903_24542# m1_12357_24542#
+ vss nfet
Xnfet$78_8 m1_2254_21786# vss m1_2384_21590# vss nfet$78
Xnfet$97_0 m1_n5351_15778# m1_n5351_15778# m1_n5461_18030# m1_n5461_18030# m1_n5225_17358#
+ vss nfet$97
Xnfet$74_73 m1_24309_25858# vss m1_21590_21786# vss nfet$74
Xnfet$74_62 m1_24188_23922# vss m1_24808_24224# vss nfet$74
Xnfet$74_51 m1_19644_25858# m1_21729_25658# m1_22522_24542# vss nfet$74
Xnfet$74_40 m1_15598_25662# m1_16442_24224# m1_17546_25658# vss nfet$74
Xnfet$83_6 m1_32193_25858# m1_32817_25662# m1_32554_23922# vss nfet$83
Xpfet$77_7 w_n11156_26804# w_n11156_26804# m1_34093_22102# m1_34843_21786# pfet$77
Xnfet$76_5 m1_649_17714# m1_649_17714# vss vss m1_6971_20470# vss nfet$76
Xpfet$91_9 w_n11156_26804# w_n11156_26804# m1_n4464_25980# m1_n4623_25487# pfet$91
Xpfet$67_28 w_n11156_26804# m1_14422_22513# m1_14422_22513# m1_13394_22102# m1_15188_21786#
+ m1_15188_21786# pfet$67
Xpfet$67_17 w_n11156_26804# m1_21456_22513# m1_21456_22513# m1_21056_22402# m1_21590_21786#
+ m1_21590_21786# pfet$67
Xnfet$74_2 m1_n7513_20152# vss m1_4509_24346# vss nfet$74
Xpfet$68_3 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_3458_19550# m1_n3218_15478#
+ m1_n3218_15478# pfet$68
Xnfet$81_3 m1_n6433_17343# vss m1_n6274_17836# vss nfet$81
Xnfet$100_5 m1_n6973_21481# m1_n6973_21481# m1_n6839_20152# m1_n6839_20152# m1_n6282_20470#
+ vss nfet$100
Xpfet$80_2 w_n11156_26804# w_n11156_26804# m1_26873_21786# pd9 pfet$80
Xpfet$66_0 w_n11156_26804# w_n11156_26804# m1_12355_15778# m1_9485_17714# pfet$66
Xpfet$73_1 w_n11156_26804# w_n11156_26804# m1_n1134_25662# m1_n1271_25858# pfet$73
Xnfet$77_73 m1_13668_17714# vss m1_16538_15778# vss nfet$77
Xnfet$77_62 m1_18665_17343# m1_20721_15778# m1_20104_16080# vss nfet$77
Xnfet$77_51 m1_n7513_20152# vss m1_22493_16080# vss nfet$77
Xnfet$77_40 m1_n2250_17343# m1_n194_15778# m1_n811_16080# vss nfet$77
Xnfet_5 m1_8692_24346# m1_8692_24346# vss vss m1_8174_24542# vss nfet
Xnfet$78_9 m1_23356_21786# vss m1_23486_21590# vss nfet$78
Xnfet$97_1 m1_n6788_16080# m1_n6788_16080# vss vss m1_n5225_17358# vss nfet$97
Xnfet$74_63 m1_14556_21786# vss m1_19644_25858# vss nfet$74
Xnfet$74_52 m1_20126_25858# vss m1_22522_24542# vss nfet$74
Xnfet$74_41 pd5 vss m1_12805_21786# vss nfet$74
Xnfet$74_30 m1_n7513_20152# vss m1_17058_24346# vss nfet$74
Xnfet$83_7 m1_32330_25662# m1_32554_23922# m1_32818_24542# vss nfet$83
Xnfet$74_74 pd8 vss m1_23356_21786# vss nfet$74
Xpfet$77_8 w_n11156_26804# m1_34093_22102# w_n11156_26804# m1_28490_22513# pfet$77
Xnfet$76_6 m1_n1133_19550# m1_n1133_19550# vss vss m1_n695_20470# vss nfet$76
Xpfet$96_0 w_n11156_26804# m1_n6380_21786# m1_n6380_21786# m1_n5019_19550# m1_n5227_20152#
+ m1_n5227_20152# pfet$96
Xpfet$67_29 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_14022_22402# m1_12805_21786#
+ m1_12805_21786# pfet$67
Xpfet$67_18 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_24573_22402# m1_23356_21786#
+ m1_23356_21786# pfet$67
Xnfet$74_3 m1_488_21786# vss m1_2912_25858# vss nfet$74
Xpfet$68_4 w_n11156_26804# m1_6107_19404# m1_6107_19404# m1_6339_19850# m1_5901_19550#
+ m1_5901_19550# pfet$68
Xnfet$81_4 m1_n7247_17714# vss m1_n4377_15778# vss nfet$81
Xnfet$100_6 m1_2590_19404# m1_2590_19404# vss vss m1_n2445_21430# vss nfet$100
Xpfet$66_1 w_n11156_26804# w_n11156_26804# m1_11381_15778# m1_11738_16080# pfet$66
Xpfet$73_2 w_n11156_26804# w_n11156_26804# m1_n1271_25858# m1_n10452_25858# pfet$73
Xnfet$77_74 m1_14482_17343# vss m1_14641_17836# vss nfet$77
Xnfet$77_63 m1_13668_17714# vss m1_14258_17518# vss nfet$77
Xnfet$77_52 m1_23007_17836# m1_24287_16080# m1_23820_18030# vss nfet$77
Xnfet$77_30 sd6 vss m1_5148_15478# vss nfet$77
Xnfet$77_41 m1_n2091_17836# m1_n1168_15778# m1_n1989_16202# vss nfet$77
Xnfet_6 m1_8076_24224# m1_8076_24224# m1_7720_24542# m1_7720_24542# m1_8174_24542#
+ vss nfet
Xnfet$97_2 m1_n6788_16080# m1_n6788_16080# m1_n7247_17714# m1_n7247_17714# m1_n6690_16398#
+ vss nfet$97
Xnfet$74_75 m1_28371_23922# vss m1_28991_24224# vss nfet$74
Xpfet$77_9 w_n11156_26804# w_n11156_26804# fout m1_34093_22102# pfet$77
Xnfet$74_64 m1_19644_25858# vss m1_19781_25662# vss nfet$74
Xnfet$74_53 m1_23827_25858# m1_24451_25662# m1_24188_23922# vss nfet$74
Xnfet$74_42 m1_15943_25858# vss m1_16085_25662# vss nfet$74
Xnfet$74_31 m1_15943_25858# vss m1_18339_24542# vss nfet$74
Xnfet$74_20 pd3 vss m1_5771_21786# vss nfet$74
Xnfet$76_7 m1_n7383_17599# m1_n7383_17599# vss vss m1_n63_20470# vss nfet$76
Xpfet$96_1 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_n5019_19550# m1_n4485_20152#
+ m1_n4485_20152# pfet$96
Xpfet$89_0 w_n11156_26804# w_n11156_26804# m1_n8625_26174# m1_n9336_24346# pfet$89
Xpfet$67_19 w_n11156_26804# m1_24973_22513# m1_24973_22513# m1_24573_22402# m1_25107_21786#
+ m1_25107_21786# pfet$67
Xnfet$107_0 m1_n927_19404# m1_n927_19404# vss vss m1_n6282_20470# vss nfet$107
Xnfet$74_4 m1_2912_25858# vss m1_3049_25662# vss nfet$74
Xpfet$68_5 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_n695_19850# m1_1103_20152#
+ m1_1103_20152# pfet$68
Xnfet$81_5 m1_n7247_17714# vss m1_n6657_17518# vss nfet$81
Xnfet$100_7 m1_6107_19404# m1_6107_19404# m1_n5227_21418# m1_n5227_21418# m1_n2445_21430#
+ vss nfet$100
Xpfet$73_3 w_n11156_26804# w_n11156_26804# m1_1607_24542# m1_n789_25858# pfet$73
Xpfet$66_2 w_n11156_26804# m1_12355_15778# m1_11738_16080# m1_10458_17836# pfet$66
Xpfet$71_0 w_n11156_26804# w_n11156_26804# m1_2384_19550# m1_n3534_17714# pfet$71
Xnfet$77_75 sd3 vss m1_17697_15478# vss nfet$77
Xnfet$77_64 m1_13668_17714# vss m1_13198_17714# vss nfet$77
Xnfet$77_53 m1_22848_17343# vss m1_23007_17836# vss nfet$77
Xnfet$77_31 m1_1933_17343# m1_3989_15778# m1_3372_16080# vss nfet$77
Xnfet$77_20 m1_1119_17714# vss m1_1709_17518# vss nfet$77
Xnfet$77_42 m1_n811_16080# vss m1_n1168_15778# vss nfet$77
Xnfet_7 m1_9180_25658# m1_9180_25658# vss vss m1_9639_25502# vss nfet
Xnfet$97_3 m1_n6172_16202# m1_n6172_16202# vss vss m1_n6690_16398# vss nfet$97
Xnfet$74_76 m1_28492_25858# vss m1_28634_25662# vss nfet$74
Xnfet$74_65 m1_28492_25858# vss m1_25107_21786# vss nfet$74
Xnfet$74_54 m1_24309_25858# vss m1_24451_25662# vss nfet$74
Xnfet$74_43 m1_15461_25858# vss m1_15598_25662# vss nfet$74
Xnfet$74_32 m1_15461_25858# m1_17546_25658# m1_18339_24542# vss nfet$74
Xnfet$74_21 m1_11278_25858# m1_11902_25662# m1_11639_23922# vss nfet$74
Xnfet$74_10 m1_7577_25858# vss m1_9973_24542# vss nfet$74
Xnfet$95_0 m1_35837_22102# vss m1_n7513_20152# vss nfet$95
Xnfet$76_8 m1_27003_19550# m1_27003_19550# vss vss m1_27441_20470# vss nfet$76
Xpfet$89_1 w_n11156_26804# m1_n8625_26174# w_n11156_26804# m1_n8848_25658# pfet$89
Xnfet$107_1 m1_n3822_20130# m1_n3822_20130# m1_n4485_20152# m1_n4485_20152# m1_n3724_20470#
+ vss nfet$107
Xnfet$74_5 m1_2912_25858# m1_3536_25662# m1_3273_23922# vss nfet$74
Xpfet$68_6 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_6339_19850# m1_8137_20152#
+ m1_8137_20152# pfet$68
Xnfet$81_6 m1_n7247_17714# vss m1_n7383_17599# vss nfet$81
Xnfet$100_8 m1_n5764_21786# m1_n5764_21786# vss vss m1_n6282_21430# vss nfet$100
Xpfet$68_30 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_24560_19550# m1_21880_15478#
+ m1_21880_15478# pfet$68
Xpfet$73_4 w_n11156_26804# w_n11156_26804# m1_488_21786# m1_n789_25858# pfet$73
Xpfet$66_3 w_n11156_26804# m1_11381_15778# m1_10560_16202# m1_10299_17343# pfet$66
Xnfet$82_10 m1_32675_25947# vss m1_35071_24542# vss nfet$82
Xpfet$71_1 w_n11156_26804# w_n11156_26804# m1_4620_20152# m1_n3218_15478# pfet$71
Xnfet$77_76 m1_14482_17343# m1_16538_15778# m1_15921_16080# vss nfet$77
Xnfet$77_65 m1_14482_17343# m1_14743_16202# m1_14258_17518# vss nfet$77
Xnfet$77_54 m1_22848_17343# m1_23109_16202# m1_22624_17518# vss nfet$77
Xnfet$77_32 m1_2092_17836# m1_3015_15778# m1_2194_16202# vss nfet$77
Xnfet$77_21 m1_1933_17343# m1_2194_16202# m1_1709_17518# vss nfet$77
Xnfet$77_10 m1_11738_16080# vss m1_11381_15778# vss nfet$77
Xnfet$77_43 sd8 vss m1_n3218_15478# vss nfet$77
Xnfet$93_20 m1_22493_16080# m1_22493_16080# m1_22034_17714# m1_22034_17714# m1_22591_16398#
+ vss nfet$93
Xnfet_8 m1_8692_24346# m1_8692_24346# m1_7577_25858# m1_7577_25858# m1_9639_25502#
+ vss nfet
Xnfet$97_4 m1_28113_15778# m1_28113_15778# m1_28003_18030# m1_28003_18030# m1_28239_17358#
+ vss nfet$97
Xnfet$74_77 m1_28010_25858# vss m1_28147_25662# vss nfet$74
Xnfet$74_66 m1_28010_25858# m1_30095_25658# m1_30888_24542# vss nfet$74
Xnfet$74_55 m1_23827_25858# vss m1_23964_25662# vss nfet$74
Xnfet$74_44 m1_15822_23922# vss m1_16442_24224# vss nfet$74
Xnfet$74_33 m1_11760_25858# vss m1_14156_24542# vss nfet$74
Xnfet$74_22 m1_11760_25858# vss m1_11902_25662# vss nfet$74
Xnfet$74_11 m1_7522_21786# vss m1_11278_25858# vss nfet$74
Xnfet$76_9 m1_25747_17714# m1_25747_17714# vss vss m1_28073_20470# vss nfet$76
Xpfet$89_2 w_n11156_26804# m1_n3651_26174# w_n11156_26804# m1_n4978_24224# pfet$89
Xnfet$88_0 m1_34843_21786# m1_34843_21786# m1_34093_22102# m1_34093_22102# m1_34329_21430#
+ vss nfet$88
Xnfet$107_2 m1_n1927_20274# m1_n1927_20274# vss vss m1_n2445_20470# vss nfet$107
Xnfet$81_7 m1_26217_17714# vss m1_26807_17518# vss nfet$81
Xnfet$74_6 m1_3049_25662# m1_3893_24224# m1_4997_25658# vss nfet$74
Xpfet$68_7 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_6975_19550# m1_965_15478#
+ m1_965_15478# pfet$68
Xpfet$94_0 w_n11156_26804# m1_n6380_21786# m1_n6380_21786# m1_n5019_19550# m1_n5227_20152#
+ m1_n5227_20152# pfet$94
Xnfet$100_9 m1_n3822_21786# m1_n3822_21786# m1_n4485_21904# m1_n4485_21904# m1_n3724_21430#
+ vss nfet$100
Xpfet$68_31 w_n11156_26804# m1_n2543_20130# m1_n2543_20130# m1_20407_19850# m1_19969_19550#
+ m1_19969_19550# pfet$68
Xpfet$68_20 w_n11156_26804# m1_n3822_21786# m1_n3822_21786# m1_14009_19550# m1_9015_17714#
+ m1_9015_17714# pfet$68
Xpfet$73_5 w_n11156_26804# w_n11156_26804# m1_326_24346# m1_n7513_20152# pfet$73
Xpfet$66_4 w_n11156_26804# m1_9485_17714# w_n11156_26804# m1_10560_16202# pfet$66
Xnfet$82_11 m1_32554_23922# vss m1_33174_24224# vss nfet$82
Xpfet$70_10 w_n11156_26804# w_n11156_26804# m1_27031_17343# m1_n10452_25858# pfet$70
Xpfet$71_2 w_n11156_26804# w_n11156_26804# m1_1103_20152# m1_n7401_15478# pfet$71
Xnfet$77_77 sd4 vss m1_13514_15478# vss nfet$77
Xnfet$77_66 m1_n7513_20152# vss m1_14127_16080# vss nfet$77
Xnfet$93_21 m1_14127_16080# m1_14127_16080# vss vss m1_15690_17358# vss nfet$93
Xnfet$77_55 m1_22034_17714# vss m1_24904_15778# vss nfet$77
Xnfet$77_44 m1_n2091_17836# m1_n811_16080# m1_n1278_18030# vss nfet$77
Xnfet$77_33 sd7 vss m1_965_15478# vss nfet$77
Xnfet$93_10 m1_1578_16080# m1_1578_16080# m1_1119_17714# m1_1119_17714# m1_1676_16398#
+ vss nfet$93
Xnfet$77_22 m1_6116_17343# m1_6377_16202# m1_5892_17518# vss nfet$77
Xnfet$77_11 m1_10299_17343# m1_12355_15778# m1_11738_16080# vss nfet$77
Xnfet_9 m1_17058_24346# m1_17058_24346# vss vss m1_16540_24542# vss nfet
Xnfet$97_5 m1_26676_16080# m1_26676_16080# vss vss m1_28239_17358# vss nfet$97
Xnfet$74_78 m1_28010_25858# m1_28634_25662# m1_28371_23922# vss nfet$74
Xnfet$74_67 m1_28492_25858# vss m1_30888_24542# vss nfet$74
Xnfet$74_56 m1_19781_25662# m1_20625_24224# m1_21729_25658# vss nfet$74
Xnfet$74_45 m1_15461_25858# m1_16085_25662# m1_15822_23922# vss nfet$74
Xnfet$74_34 m1_11278_25858# m1_13363_25658# m1_14156_24542# vss nfet$74
Xnfet$74_23 m1_11278_25858# vss m1_11415_25662# vss nfet$74
Xnfet$74_12 m1_7577_25858# vss m1_7522_21786# vss nfet$74
Xnfet$88_1 m1_28490_22513# m1_28490_22513# vss vss m1_34329_21430# vss nfet$88
Xpfet$89_3 w_n11156_26804# w_n11156_26804# m1_n3651_26174# m1_n3541_23922# pfet$89
Xnfet$107_3 m1_n2543_20130# m1_n2543_20130# m1_n5227_20152# m1_n5227_20152# m1_n2445_20470#
+ vss nfet$107
Xpfet$73_10 w_n11156_26804# w_n11156_26804# m1_35071_24542# m1_32675_25947# pfet$73
Xnfet$81_8 m1_n7513_20152# vss m1_26676_16080# vss nfet$81
Xnfet$74_7 m1_3049_25662# m1_3273_23922# m1_3537_24542# vss nfet$74
Xpfet$68_8 w_n11156_26804# m1_9624_19404# m1_9624_19404# m1_10492_19550# m1_4832_17714#
+ m1_4832_17714# pfet$68
Xpfet$94_1 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_n5019_19550# m1_n4485_20152#
+ m1_n4485_20152# pfet$94
Xpfet$87_0 w_n11156_26804# m1_n10309_25662# m1_n10572_23922# m1_n10796_25662# pfet$87
Xnfet$105_0 m1_n8283_20611# vss m1_n8283_19850# vss nfet$105
Xpfet$68_32 w_n11156_26804# m1_n2543_20130# m1_n2543_20130# m1_21043_19550# m1_17381_17714#
+ m1_17381_17714# pfet$68
Xpfet$68_21 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_13373_19850# m1_15171_20152#
+ m1_15171_20152# pfet$68
Xpfet$73_6 w_n11156_26804# w_n11156_26804# m1_n290_24224# m1_n910_23922# pfet$73
Xpfet$66_5 w_n11156_26804# m1_7198_15778# m1_6377_16202# m1_6116_17343# pfet$66
Xpfet$68_10 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_9856_19850# m1_11654_20152#
+ m1_11654_20152# pfet$68
Xnfet$82_12 m1_32675_25947# vss m1_28624_21786# vss nfet$82
Xpfet$70_11 w_n11156_26804# w_n11156_26804# m1_26807_17518# m1_26217_17714# pfet$70
Xpfet$71_3 w_n11156_26804# w_n11156_26804# m1_5901_19550# m1_649_17714# pfet$71
Xnfet$77_78 m1_14641_17836# m1_15564_15778# m1_14743_16202# vss nfet$77
Xnfet$93_22 m1_15564_15778# m1_15564_15778# m1_15454_18030# m1_15454_18030# m1_15690_17358#
+ vss nfet$93
Xnfet$77_67 m1_17381_17714# vss m1_14482_17343# vss nfet$77
Xnfet$77_56 m1_24287_16080# vss m1_23930_15778# vss nfet$77
Xnfet$77_45 m1_n3064_17714# vss m1_n194_15778# vss nfet$77
Xnfet$77_34 m1_n2250_17343# vss m1_n2091_17836# vss nfet$77
Xnfet$77_23 m1_5302_17714# vss m1_4832_17714# vss nfet$77
Xnfet$77_12 m1_9485_17714# vss m1_12355_15778# vss nfet$77
Xnfet$93_11 m1_6377_16202# m1_6377_16202# vss vss m1_5859_16398# vss nfet$93
Xnfet$97_6 m1_27292_16202# m1_27292_16202# vss vss m1_26774_16398# vss nfet$97
Xnfet$74_68 m1_n7513_20152# vss m1_29607_24346# vss nfet$74
Xnfet$74_57 m1_20126_25858# vss m1_20268_25662# vss nfet$74
Xnfet$74_46 m1_20126_25858# vss m1_18073_21786# vss nfet$74
Xnfet$74_35 m1_15598_25662# m1_15822_23922# m1_16086_24542# vss nfet$74
Xnfet$74_24 m1_7095_25858# m1_7719_25662# m1_7456_23922# vss nfet$74
Xnfet$74_13 m1_11415_25662# m1_11639_23922# m1_11903_24542# vss nfet$74
Xnfet$74_79 pd7 vss m1_19839_21786# vss nfet$74
Xnfet$88_2 m1_9645_21447# m1_9645_21447# vss vss m1_30492_21430# vss nfet$88
Xpfet$89_4 w_n11156_26804# m1_n10452_25858# w_n11156_26804# m1_n4362_24346# pfet$89
Xnfet$107_4 m1_n3206_20274# m1_n3206_20274# vss vss m1_n3724_20470# vss nfet$107
Xpfet$73_11 w_n11156_26804# w_n11156_26804# m1_32817_25662# m1_32675_25947# pfet$73
Xnfet$81_9 m1_n10452_25858# vss m1_27031_17343# vss nfet$81
Xnfet$74_8 m1_3394_25858# vss m1_3536_25662# vss nfet$74
Xpfet$68_9 w_n11156_26804# m1_9624_19404# m1_9624_19404# m1_9856_19850# m1_9418_19550#
+ m1_9418_19550# pfet$68
Xpfet$94_2 w_n11156_26804# m1_n5764_21786# m1_n5764_21786# m1_n5019_22344# m1_n5227_21418#
+ m1_n5227_21418# pfet$94
Xpfet$87_1 w_n11156_26804# m1_n9952_24224# m1_n8848_25658# m1_n10933_25858# pfet$87
Xnfet$93_0 m1_7198_15778# m1_7198_15778# m1_7088_18030# m1_7088_18030# m1_7324_17358#
+ vss nfet$93
Xnfet$105_1 m1_n7513_20152# m1_n8283_19850# vss vss nfet$105
Xpfet$73_7 w_n11156_26804# w_n11156_26804# m1_32330_25662# m1_32193_25858# pfet$73
Xpfet$68_33 w_n11156_26804# m1_n3206_20274# m1_n3206_20274# m1_24560_19550# m1_21564_17714#
+ m1_21564_17714# pfet$68
Xpfet$68_22 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_14009_19550# m1_9331_15478#
+ m1_9331_15478# pfet$68
Xpfet$66_6 w_n11156_26804# w_n11156_26804# m1_7198_15778# m1_7555_16080# pfet$66
Xpfet$68_11 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_10492_19550# m1_5148_15478#
+ m1_5148_15478# pfet$68
Xnfet$82_13 m1_32675_25947# vss m1_32817_25662# vss nfet$82
Xpfet$70_12 w_n11156_26804# w_n11156_26804# m1_26676_16080# m1_n7513_20152# pfet$70
Xpfet$71_4 w_n11156_26804# w_n11156_26804# m1_12935_19550# m1_9015_17714# pfet$71
Xnfet$77_79 m1_15921_16080# vss m1_15564_15778# vss nfet$77
Xnfet$93_23 m1_18926_16202# m1_18926_16202# vss vss m1_18408_16398# vss nfet$93
Xnfet$77_68 m1_18665_17343# m1_18926_16202# m1_18441_17518# vss nfet$77
Xnfet$77_57 m1_22848_17343# m1_24904_15778# m1_24287_16080# vss nfet$77
Xnfet$77_46 m1_22034_17714# vss m1_21564_17714# vss nfet$77
Xnfet$77_24 m1_4832_17714# vss m1_1933_17343# vss nfet$77
Xnfet$77_13 m1_10458_17836# m1_11381_15778# m1_10560_16202# vss nfet$77
Xnfet$77_35 m1_n7513_20152# vss m1_5761_16080# vss nfet$77
Xnfet$93_12 m1_n1168_15778# m1_n1168_15778# m1_n1278_18030# m1_n1278_18030# m1_n1042_17358#
+ vss nfet$93
Xnfet$97_7 m1_26676_16080# m1_26676_16080# m1_26217_17714# m1_26217_17714# m1_26774_16398#
+ vss nfet$97
Xnfet$74_69 m1_24309_25858# vss m1_26705_24542# vss nfet$74
Xnfet$74_58 m1_20005_23922# vss m1_20625_24224# vss nfet$74
Xnfet$74_47 m1_23964_25662# m1_24188_23922# m1_24452_24542# vss nfet$74
Xnfet$74_36 m1_11760_25858# vss m1_11039_21786# vss nfet$74
Xnfet$74_25 m1_7232_25662# m1_8076_24224# m1_9180_25658# vss nfet$74
Xnfet$74_14 m1_n7513_20152# vss m1_8692_24346# vss nfet$74
Xnfet$88_3 m1_7388_22513# m1_7388_22513# m1_30256_22102# m1_30256_22102# m1_30492_21430#
+ vss nfet$88
Xpfet$89_5 w_n11156_26804# w_n11156_26804# m1_n10308_24542# m1_n9952_24224# pfet$89
Xnfet$107_5 m1_n6973_21481# m1_n6973_21481# m1_n6839_20152# m1_n6839_20152# m1_n6282_20470#
+ vss nfet$107
Xpfet$73_12 w_n11156_26804# w_n11156_26804# m1_32193_25858# m1_25107_21786# pfet$73
Xnfet$74_9 m1_3273_23922# vss m1_3893_24224# vss nfet$74
Xnfet$93_1 m1_5761_16080# m1_5761_16080# vss vss m1_7324_17358# vss nfet$93
Xpfet$94_3 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_n5019_22344# m1_n4485_21904#
+ m1_n4485_21904# pfet$94
Xpfet$87_2 w_n11156_26804# m1_n4362_24346# m1_n4847_25662# m1_n4464_25980# pfet$87
Xnfet$86_0 m1_11039_21786# m1_11039_21786# vss vss m1_9877_21586# vss nfet$86
Xpfet$73_8 w_n11156_26804# w_n11156_26804# m1_33174_24224# m1_32554_23922# pfet$73
Xpfet$68_34 w_n11156_26804# m1_n3206_20274# m1_n3206_20274# m1_23924_19850# m1_23486_19550#
+ m1_23486_19550# pfet$68
Xpfet$68_23 w_n11156_26804# w_n11156_26804# w_n11156_26804# m1_16890_19850# m1_18688_20152#
+ m1_18688_20152# pfet$68
Xpfet$68_12 w_n11156_26804# m1_6107_19404# m1_6107_19404# m1_6975_19550# m1_649_17714#
+ m1_649_17714# pfet$68
Xnfet$105_2 m1_n8145_21908# vss m1_n8283_20611# vss nfet$105
Xpfet$66_7 w_n11156_26804# w_n11156_26804# m1_6275_17836# m1_6116_17343# pfet$66
Xpfet$92_0 w_n11156_26804# w_n11156_26804# m1_n7186_25858# m1_n10452_25858# pfet$92
Xpfet$70_13 w_n11156_26804# w_n11156_26804# m1_25747_17714# m1_26217_17714# pfet$70
Xpfet$71_5 w_n11156_26804# w_n11156_26804# m1_8137_20152# m1_965_15478# pfet$71
Xnfet$93_24 m1_18310_16080# m1_18310_16080# m1_17851_17714# m1_17851_17714# m1_18408_16398#
+ vss nfet$93
Xnfet$77_69 m1_17851_17714# vss m1_17381_17714# vss nfet$77
Xnfet$77_58 m1_23007_17836# m1_23930_15778# m1_23109_16202# vss nfet$77
Xnfet$77_47 m1_22034_17714# vss m1_22624_17518# vss nfet$77
Xnfet$77_25 m1_2092_17836# m1_3372_16080# m1_2905_18030# vss nfet$77
Xnfet$77_14 m1_6116_17343# m1_8172_15778# m1_7555_16080# vss nfet$77
Xnfet$77_36 m1_n3064_17714# vss m1_n2474_17518# vss nfet$77
Xnfet$93_13 m1_n2605_16080# m1_n2605_16080# vss vss m1_n1042_17358# vss nfet$93
Xnfet$74_59 m1_19644_25858# m1_20268_25662# m1_20005_23922# vss nfet$74
Xnfet$74_48 m1_18073_21786# vss m1_23827_25858# vss nfet$74
Xnfet$74_37 m1_11039_21786# vss m1_15461_25858# vss nfet$74
Xnfet$74_26 m1_7095_25858# m1_9180_25658# m1_9973_24542# vss nfet$74
Xnfet$74_15 m1_7232_25662# m1_7456_23922# m1_7720_24542# vss nfet$74
Xnfet$88_4 m1_3871_22513# m1_3871_22513# vss vss m1_31771_21430# vss nfet$88
Xpfet$89_6 w_n11156_26804# m1_n10308_24542# w_n11156_26804# m1_n9336_24346# pfet$89
Xpfet$73_13 w_n11156_26804# w_n11156_26804# m1_33790_24346# m1_n7513_20152# pfet$73
Xnfet$79_0 m1_n3534_17714# vss m1_2384_19550# vss nfet$79
Xnfet$93_2 m1_9944_16080# m1_9944_16080# vss vss m1_11507_17358# vss nfet$93
Xpfet$87_3 w_n11156_26804# m1_n3184_24224# m1_n3651_26174# m1_n4623_25487# pfet$87
Xnfet$86_1 m1_11671_21786# m1_11671_21786# vss vss m1_10509_21586# vss nfet$86
Xpfet$68_13 w_n11156_26804# m1_n927_19404# m1_n927_19404# m1_n695_19850# m1_n1133_19550#
+ m1_n1133_19550# pfet$68
Xnfet$105_3 m1_n8283_19850# m1_n8283_20611# vss vss nfet$105
Xpfet$68_35 w_n11156_26804# m1_n3822_21786# m1_n3822_21786# m1_13373_19850# m1_12935_19550#
+ m1_12935_19550# pfet$68
Xpfet$73_9 w_n11156_26804# w_n11156_26804# m1_28624_21786# m1_32675_25947# pfet$73
Xpfet$68_24 w_n11156_26804# m1_n1927_20274# m1_n1927_20274# m1_16890_19850# m1_16452_19550#
+ m1_16452_19550# pfet$68
Xpfet$66_8 w_n11156_26804# w_n11156_26804# m1_9331_15478# sd5 pfet$66
Xpfet$92_1 w_n11156_26804# m1_n7186_25858# w_n11156_26804# m1_n6111_25858# pfet$92
Xpfet$85_0 w_n11156_26804# w_n11156_26804# m1_n7513_20152# m1_35837_22102# pfet$85
Xnfet$103_0 m1_n10933_25858# m1_n8848_25658# m1_n8055_24542# vss nfet$103
Xpfet$71_6 w_n11156_26804# w_n11156_26804# m1_9418_19550# m1_4832_17714# pfet$71
Xnfet$77_59 m1_17851_17714# vss m1_20721_15778# vss nfet$77
Xnfet$77_48 m1_18824_17836# m1_20104_16080# m1_19637_18030# vss nfet$77
Xnfet$77_26 m1_5302_17714# vss m1_5892_17518# vss nfet$77
Xnfet$77_15 m1_5302_17714# vss m1_8172_15778# vss nfet$77
Xnfet$77_37 m1_n7513_20152# vss m1_n2605_16080# vss nfet$77
Xnfet$93_25 m1_14743_16202# m1_14743_16202# vss vss m1_14225_16398# vss nfet$93
Xnfet$93_14 m1_n2605_16080# m1_n2605_16080# m1_n3064_17714# m1_n3064_17714# m1_n2507_16398#
+ vss nfet$93
Xpfet_90 w_n11156_26804# w_n11156_26804# m1_24309_25858# m1_25424_24346# pfet
Xnfet$74_49 m1_19781_25662# m1_20005_23922# m1_20269_24542# vss nfet$74
Xnfet$74_38 m1_n7513_20152# vss m1_12875_24346# vss nfet$74
Xpfet$66_90 w_n11156_26804# m1_19747_15778# m1_18926_16202# m1_18665_17343# pfet$66
Xnfet$74_27 m1_7577_25858# vss m1_7719_25662# vss nfet$74
Xnfet$74_16 m1_4005_21786# vss m1_7095_25858# vss nfet$74
Xpfet$89_7 w_n11156_26804# w_n11156_26804# m1_n10452_25858# m1_n4978_24224# pfet$89
Xnfet$88_5 m1_354_22513# m1_354_22513# m1_31535_22102# m1_31535_22102# m1_31771_21430#
+ vss nfet$88
.ends

.subckt pfet$4 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$2 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$3 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt nfet$1 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$3 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$1 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$4 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$2 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt asc_drive_buffer vss in vdd out
Xpfet$4_0 vdd vdd m1_3466_n454# in pfet$4
Xpfet$2_0 m1_4274_n1060# vdd vdd m1_4274_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ vdd m1_4002_n1060# m1_4002_n1060# pfet$2
Xnfet$3_0 m1_3466_n454# vss m1_4002_n1060# vss nfet$3
Xnfet$1_0 m1_4274_n1060# vss m1_4002_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ m1_4274_n1060# vss m1_4002_n1060# vss nfet$1
Xpfet$3_0 vdd vdd m1_4002_n1060# m1_3466_n454# pfet$3
Xpfet$1_0 out out m1_4274_n1060# vdd m1_4274_n1060# out vdd vdd m1_4274_n1060# out
+ m1_4274_n1060# m1_4274_n1060# out m1_4274_n1060# vdd m1_4274_n1060# vdd m1_4274_n1060#
+ pfet$1
Xnfet$4_0 in vss m1_3466_n454# vss nfet$4
Xnfet$2_0 out out vss m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# m1_4274_n1060#
+ m1_4274_n1060# out m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# vss vss
+ nfet$2
.ends

.subckt pfet$30 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$29 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$28 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$27 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$26 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$30 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$29 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$28 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$27 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$26 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt asc_hysteresis_buffer vss in vdd out
Xpfet$30_0 vdd vdd m1_884_42# m1_1156_42# pfet$30
Xnfet$29_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$29
Xpfet$28_0 vdd vdd m1_348_648# in pfet$28
Xnfet$27_0 m1_348_648# vss m1_884_42# vss nfet$27
Xpfet$26_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd m1_884_42#
+ m1_884_42# pfet$26
Xnfet$30_0 m1_1156_42# vss m1_884_42# vss nfet$30
Xpfet$29_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$29
Xnfet$28_0 in vss m1_348_648# vss nfet$28
Xpfet$27_0 vdd vdd m1_884_42# m1_348_648# pfet$27
Xnfet$26_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$26
.ends

.subckt nfet$17 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$8 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$16 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$15 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$6 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$9 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$14 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$13 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$7 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$12 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$11 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$5 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$10 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$19 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$18 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$9 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$17 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$16 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$7 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$15 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$14 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$5 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$8 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$13 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$12 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$6 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$11 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$10 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$19 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$18 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt asc_lock_detector_20250826 ref vdd div lock vss
Xnfet$17_0 m1_n4030_5270# vss m1_n2336_5099# vss nfet$17
Xpfet$8_0 m1_7448_n340# vdd vdd m1_7448_n340# m1_7176_n340# m1_7176_n340# m1_7448_n340#
+ vdd m1_7176_n340# m1_7176_n340# pfet$8
Xpfet$16_0 vdd vdd vdd m1_n3798_6028# div div pfet$16
Xpfet$8_1 m1_11642_n340# vdd vdd m1_11642_n340# m1_11370_n340# m1_11370_n340# m1_11642_n340#
+ vdd m1_11370_n340# m1_11370_n340# pfet$8
Xpfet$16_1 vdd m1_n4030_5270# m1_n4030_5270# m1_n3798_6028# m1_n6066_7868# m1_n6066_7868#
+ pfet$16
Xpfet$8_2 m1_3254_n340# vdd vdd m1_3254_n340# m1_2982_n340# m1_2982_n340# m1_3254_n340#
+ vdd m1_2982_n340# m1_2982_n340# pfet$8
Xnfet$15_0 m1_n14454_7868# vss m1_n12216_5099# vss nfet$15
Xpfet$8_3 m1_n940_n340# vdd vdd m1_n940_n340# m1_n1212_n340# m1_n1212_n340# m1_n940_n340#
+ vdd m1_n1212_n340# m1_n1212_n340# pfet$8
Xpfet$6_0 vdd vdd m1_7176_n340# m1_6640_1478# pfet$6
Xnfet$9_0 m1_n8022_5099# vss m1_n7486_4493# vss nfet$9
Xnfet$15_1 div vss m1_n16410_5099# vss nfet$15
Xpfet$14_0 vdd vdd m1_n11680_4493# m1_n12216_5099# pfet$14
Xpfet$8_4 m1_n940_4493# vdd vdd m1_n940_4493# m1_n1212_4493# m1_n1212_4493# m1_n940_4493#
+ vdd m1_n1212_4493# m1_n1212_4493# pfet$8
Xpfet$6_1 vdd vdd m1_11370_n340# m1_10834_1478# pfet$6
Xnfet$9_1 m1_n16410_5099# vss m1_n15874_4493# vss nfet$9
Xnfet$15_2 m1_n10260_7868# vss m1_n8022_5099# vss nfet$15
Xpfet$14_1 vdd vdd m1_n7486_4493# m1_n8022_5099# pfet$14
Xpfet$8_5 m1_11642_4493# vdd vdd m1_11642_4493# m1_11370_4493# m1_11370_4493# m1_11642_4493#
+ vdd m1_11370_4493# m1_11370_4493# pfet$8
Xpfet$6_2 vdd vdd m1_2982_n340# m1_2446_1478# pfet$6
Xnfet$9_2 m1_n12216_5099# vss m1_n11680_4493# vss nfet$9
Xpfet$8_6 m1_3254_4493# vdd vdd m1_3254_4493# m1_2982_4493# m1_2982_4493# m1_3254_4493#
+ vdd m1_2982_4493# m1_2982_4493# pfet$8
Xnfet$13_0 m1_17215_2028# m1_17215_2028# m1_17926_34# m1_17926_34# m1_18162_712# vss
+ nfet$13
Xpfet$14_2 vdd vdd m1_n15874_4493# m1_n16410_5099# pfet$14
Xpfet$6_3 vdd vdd m1_n1212_n340# m1_n1748_1478# pfet$6
Xnfet$13_1 m1_17703_788# m1_17703_788# vss vss m1_18162_712# vss nfet$13
Xnfet$7_0 m1_3254_n340# vss m1_2982_n340# m1_2982_n340# m1_2982_n340# m1_3254_n340#
+ m1_3254_n340# vss m1_2982_n340# vss nfet$7
Xpfet$8_7 m1_7448_4493# vdd vdd m1_7448_4493# m1_7176_4493# m1_7176_4493# m1_7448_4493#
+ vdd m1_7176_4493# m1_7176_4493# pfet$8
Xpfet$12_0 m1_n10260_7868# m1_n10260_7868# m1_n11408_4493# vdd m1_n11408_4493# m1_n10260_7868#
+ vdd vdd m1_n11408_4493# m1_n10260_7868# m1_n11408_4493# m1_n11408_4493# m1_n10260_7868#
+ m1_n11408_4493# vdd m1_n11408_4493# vdd m1_n11408_4493# pfet$12
Xpfet$6_4 vdd vdd m1_n1212_4493# m1_n1748_5099# pfet$6
Xnfet$7_1 m1_7448_n340# vss m1_7176_n340# m1_7176_n340# m1_7176_n340# m1_7448_n340#
+ m1_7448_n340# vss m1_7176_n340# vss nfet$7
Xnfet$13_2 m1_16599_2028# m1_16599_2028# m1_16243_1828# m1_16243_1828# m1_16697_1672#
+ vss nfet$13
Xpfet$12_1 m1_n6066_7868# m1_n6066_7868# m1_n7214_4493# vdd m1_n7214_4493# m1_n6066_7868#
+ vdd vdd m1_n7214_4493# m1_n6066_7868# m1_n7214_4493# m1_n7214_4493# m1_n6066_7868#
+ m1_n7214_4493# vdd m1_n7214_4493# vdd m1_n7214_4493# pfet$12
Xpfet$6_5 vdd vdd m1_2982_4493# m1_2446_5099# pfet$6
Xnfet$13_3 m1_17215_2028# m1_17215_2028# vss vss m1_16697_1672# vss nfet$13
Xnfet$7_2 m1_11642_n340# vss m1_11370_n340# m1_11370_n340# m1_11370_n340# m1_11642_n340#
+ m1_11642_n340# vss m1_11370_n340# vss nfet$7
Xpfet$6_6 vdd vdd m1_7176_4493# m1_6640_5099# pfet$6
Xnfet$11_0 m1_8596_n340# vss m1_10834_1478# vss nfet$11
Xpfet$12_2 m1_n14454_7868# m1_n14454_7868# m1_n15602_4493# vdd m1_n15602_4493# m1_n14454_7868#
+ vdd vdd m1_n15602_4493# m1_n14454_7868# m1_n15602_4493# m1_n15602_4493# m1_n14454_7868#
+ m1_n15602_4493# vdd m1_n15602_4493# vdd m1_n15602_4493# pfet$12
Xnfet$7_3 m1_n940_n340# vss m1_n1212_n340# m1_n1212_n340# m1_n1212_n340# m1_n940_n340#
+ m1_n940_n340# vss m1_n1212_n340# vss nfet$7
Xnfet$5_0 m1_8596_n340# m1_8596_n340# vss m1_7448_n340# m1_7448_n340# m1_8596_n340#
+ vss m1_7448_n340# m1_7448_n340# m1_7448_n340# m1_8596_n340# m1_7448_n340# m1_7448_n340#
+ m1_8596_n340# vss m1_7448_n340# vss vss nfet$5
Xnfet$11_1 m1_4402_n340# vss m1_6640_1478# vss nfet$11
Xnfet$13_4 m1_17215_5644# m1_17215_5644# vss vss m1_16697_5840# vss nfet$13
Xpfet$6_7 vdd vdd m1_11370_4493# m1_10834_5099# pfet$6
Xpfet$10_0 vdd m1_16599_2028# m1_17703_788# m1_15618_394# pfet$10
Xnfet$7_4 m1_11642_4493# vss m1_11370_4493# m1_11370_4493# m1_11370_4493# m1_11642_4493#
+ m1_11642_4493# vss m1_11370_4493# vss nfet$7
Xnfet$13_5 m1_16599_5522# m1_16599_5522# m1_16243_5840# m1_16243_5840# m1_16697_5840#
+ vss nfet$13
Xnfet$5_1 m1_4402_n340# m1_4402_n340# vss m1_3254_n340# m1_3254_n340# m1_4402_n340#
+ vss m1_3254_n340# m1_3254_n340# m1_3254_n340# m1_4402_n340# m1_3254_n340# m1_3254_n340#
+ m1_4402_n340# vss m1_3254_n340# vss vss nfet$5
Xnfet$11_2 ref vss m1_n1748_1478# vss nfet$11
Xpfet$10_1 vdd m1_16242_n208# m1_15979_2344# m1_15755_n208# pfet$10
Xnfet$7_5 m1_7448_4493# vss m1_7176_4493# m1_7176_4493# m1_7176_4493# m1_7448_4493#
+ m1_7448_4493# vss m1_7176_4493# vss nfet$7
Xnfet$13_6 m1_17215_5644# m1_17215_5644# m1_17926_7472# m1_17926_7472# m1_18162_6800#
+ vss nfet$13
Xnfet$5_2 m1_12790_n340# m1_12790_n340# vss m1_11642_n340# m1_11642_n340# m1_12790_n340#
+ vss m1_11642_n340# m1_11642_n340# m1_11642_n340# m1_12790_n340# m1_11642_n340# m1_11642_n340#
+ m1_12790_n340# vss m1_11642_n340# vss vss nfet$5
Xpfet$10_2 vdd m1_15979_2344# m1_16243_1828# m1_15618_394# pfet$10
Xnfet$11_3 m1_n2336_5099# vss m1_n1748_5099# vss nfet$11
Xnfet$7_6 m1_n940_4493# vss m1_n1212_4493# m1_n1212_4493# m1_n1212_4493# m1_n940_4493#
+ m1_n940_4493# vss m1_n1212_4493# vss nfet$7
Xnfet$13_7 m1_17703_6956# m1_17703_6956# vss vss m1_18162_6800# vss nfet$13
Xnfet$11_4 m1_8596_7868# vss m1_10834_5099# vss nfet$11
Xnfet$5_3 m1_208_n340# m1_208_n340# vss m1_n940_n340# m1_n940_n340# m1_208_n340# vss
+ m1_n940_n340# m1_n940_n340# m1_n940_n340# m1_208_n340# m1_n940_n340# m1_n940_n340#
+ m1_208_n340# vss m1_n940_n340# vss vss nfet$5
Xpfet$10_3 vdd m1_17703_788# m1_18496_1828# m1_15755_n208# pfet$10
Xnfet$7_7 m1_3254_4493# vss m1_2982_4493# m1_2982_4493# m1_2982_4493# m1_3254_4493#
+ m1_3254_4493# vss m1_2982_4493# vss nfet$7
Xnfet$5_4 m1_12790_7868# m1_12790_7868# vss m1_11642_4493# m1_11642_4493# m1_12790_7868#
+ vss m1_11642_4493# m1_11642_4493# m1_11642_4493# m1_12790_7868# m1_11642_4493# m1_11642_4493#
+ m1_12790_7868# vss m1_11642_4493# vss vss nfet$5
Xpfet$19_0 vdd vdd lock m1_19675_2344# pfet$19
Xnfet$11_5 m1_4402_7868# vss m1_6640_5099# vss nfet$11
Xpfet$10_4 vdd m1_17703_6956# m1_18496_5840# m1_15755_6960# pfet$10
Xnfet$5_5 m1_8596_7868# m1_8596_7868# vss m1_7448_4493# m1_7448_4493# m1_8596_7868#
+ vss m1_7448_4493# m1_7448_4493# m1_7448_4493# m1_8596_7868# m1_7448_4493# m1_7448_4493#
+ m1_8596_7868# vss m1_7448_4493# vss vss nfet$5
Xnfet$11_6 m1_208_n340# vss m1_2446_1478# vss nfet$11
Xpfet$10_5 vdd m1_15979_5220# m1_16243_5840# m1_15618_7156# pfet$10
Xnfet$5_6 m1_208_7868# m1_208_7868# vss m1_n940_4493# m1_n940_4493# m1_208_7868# vss
+ m1_n940_4493# m1_n940_4493# m1_n940_4493# m1_208_7868# m1_n940_4493# m1_n940_4493#
+ m1_208_7868# vss m1_n940_4493# vss vss nfet$5
Xnfet$18_0 m1_19469_4920# m1_19469_4920# m1_19675_2344# m1_19675_2344# m1_19911_1672#
+ vss nfet$18
Xnfet$11_7 m1_208_7868# vss m1_2446_5099# vss nfet$11
Xpfet$10_6 vdd m1_16599_5522# m1_17703_6956# m1_15618_7156# pfet$10
Xpfet$9_0 vdd vdd m1_16599_2028# m1_15979_2344# pfet$9
Xnfet$5_7 m1_4402_7868# m1_4402_7868# vss m1_3254_4493# m1_3254_4493# m1_4402_7868#
+ vss m1_3254_4493# m1_3254_4493# m1_3254_4493# m1_4402_7868# m1_3254_4493# m1_3254_4493#
+ m1_4402_7868# vss m1_3254_4493# vss vss nfet$5
Xnfet$18_1 m1_19469_1832# m1_19469_1832# vss vss m1_19911_1672# vss nfet$18
Xpfet$17_0 vdd vdd m1_n2336_5099# m1_n4030_5270# pfet$17
Xpfet$10_7 vdd m1_16242_6960# m1_15979_5220# m1_15755_6960# pfet$10
Xpfet$9_1 vdd vdd m1_16242_n208# m1_n2336_5099# pfet$9
Xpfet$9_2 vdd vdd m1_15755_n208# m1_15618_394# pfet$9
Xnfet$16_0 div m1_n4030_5270# vss vss nfet$16
Xpfet$9_3 vdd vdd m1_18496_1828# m1_17926_34# pfet$9
Xpfet$7_0 m1_8596_n340# m1_8596_n340# m1_7448_n340# vdd m1_7448_n340# m1_8596_n340#
+ vdd vdd m1_7448_n340# m1_8596_n340# m1_7448_n340# m1_7448_n340# m1_8596_n340# m1_7448_n340#
+ vdd m1_7448_n340# vdd m1_7448_n340# pfet$7
Xnfet$16_1 m1_n6066_7868# vss m1_n4030_5270# vss nfet$16
Xpfet$9_4 vdd vdd m1_15618_394# m1_12790_n340# pfet$9
Xpfet$15_0 vdd vdd m1_n8022_5099# m1_n10260_7868# pfet$15
Xpfet$7_1 m1_12790_n340# m1_12790_n340# m1_11642_n340# vdd m1_11642_n340# m1_12790_n340#
+ vdd vdd m1_11642_n340# m1_12790_n340# m1_11642_n340# m1_11642_n340# m1_12790_n340#
+ m1_11642_n340# vdd m1_11642_n340# vdd m1_11642_n340# pfet$7
Xpfet$15_1 vdd vdd m1_n16410_5099# div pfet$15
Xpfet$9_5 vdd vdd m1_17215_2028# vss pfet$9
Xpfet$7_2 m1_4402_n340# m1_4402_n340# m1_3254_n340# vdd m1_3254_n340# m1_4402_n340#
+ vdd vdd m1_3254_n340# m1_4402_n340# m1_3254_n340# m1_3254_n340# m1_4402_n340# m1_3254_n340#
+ vdd m1_3254_n340# vdd m1_3254_n340# pfet$7
Xnfet$14_0 m1_15979_2344# vss m1_16599_2028# vss nfet$14
Xpfet$9_6 vdd vdd m1_19469_1832# m1_17926_34# pfet$9
Xpfet$15_2 vdd vdd m1_n12216_5099# m1_n14454_7868# pfet$15
Xnfet$14_10 m1_12790_7868# vss m1_15618_7156# vss nfet$14
Xpfet$7_3 m1_208_n340# m1_208_n340# m1_n940_n340# vdd m1_n940_n340# m1_208_n340# vdd
+ vdd m1_n940_n340# m1_208_n340# m1_n940_n340# m1_n940_n340# m1_208_n340# m1_n940_n340#
+ vdd m1_n940_n340# vdd m1_n940_n340# pfet$7
Xpfet$5_0 vdd vdd m1_6640_1478# m1_4402_n340# pfet$5
Xnfet$8_0 m1_n6066_7868# m1_n6066_7868# vss m1_n7214_4493# m1_n7214_4493# m1_n6066_7868#
+ vss m1_n7214_4493# m1_n7214_4493# m1_n7214_4493# m1_n6066_7868# m1_n7214_4493# m1_n7214_4493#
+ m1_n6066_7868# vss m1_n7214_4493# vss vss nfet$8
Xnfet$14_1 m1_15618_394# vss m1_15755_n208# vss nfet$14
Xpfet$13_0 m1_n11408_4493# vdd vdd m1_n11408_4493# m1_n11680_4493# m1_n11680_4493#
+ m1_n11408_4493# vdd m1_n11680_4493# m1_n11680_4493# pfet$13
Xpfet$9_7 vdd vdd m1_17215_5644# vss pfet$9
Xnfet$14_11 m1_15979_5220# vss m1_16599_5522# vss nfet$14
Xpfet$5_1 vdd vdd m1_10834_1478# m1_8596_n340# pfet$5
Xpfet$7_4 m1_208_7868# m1_208_7868# m1_n940_4493# vdd m1_n940_4493# m1_208_7868# vdd
+ vdd m1_n940_4493# m1_208_7868# m1_n940_4493# m1_n940_4493# m1_208_7868# m1_n940_4493#
+ vdd m1_n940_4493# vdd m1_n940_4493# pfet$7
Xnfet$8_1 m1_n14454_7868# m1_n14454_7868# vss m1_n15602_4493# m1_n15602_4493# m1_n14454_7868#
+ vss m1_n15602_4493# m1_n15602_4493# m1_n15602_4493# m1_n14454_7868# m1_n15602_4493#
+ m1_n15602_4493# m1_n14454_7868# vss m1_n15602_4493# vss vss nfet$8
Xnfet$14_2 m1_n2336_5099# vss m1_16242_n208# vss nfet$14
Xnfet$14_12 m1_15618_7156# vss m1_15755_6960# vss nfet$14
Xpfet$7_5 m1_12790_7868# m1_12790_7868# m1_11642_4493# vdd m1_11642_4493# m1_12790_7868#
+ vdd vdd m1_11642_4493# m1_12790_7868# m1_11642_4493# m1_11642_4493# m1_12790_7868#
+ m1_11642_4493# vdd m1_11642_4493# vdd m1_11642_4493# pfet$7
Xpfet$9_8 vdd vdd m1_19469_4920# m1_17926_7472# pfet$9
Xpfet$13_1 m1_n7214_4493# vdd vdd m1_n7214_4493# m1_n7486_4493# m1_n7486_4493# m1_n7214_4493#
+ vdd m1_n7486_4493# m1_n7486_4493# pfet$13
Xpfet$5_2 vdd vdd m1_n1748_1478# ref pfet$5
Xnfet$8_2 m1_n10260_7868# m1_n10260_7868# vss m1_n11408_4493# m1_n11408_4493# m1_n10260_7868#
+ vss m1_n11408_4493# m1_n11408_4493# m1_n11408_4493# m1_n10260_7868# m1_n11408_4493#
+ m1_n11408_4493# m1_n10260_7868# vss m1_n11408_4493# vss vss nfet$8
Xpfet$9_10 vdd vdd m1_15618_7156# m1_12790_7868# pfet$9
Xpfet$9_9 vdd vdd m1_18496_5840# m1_17926_7472# pfet$9
Xnfet$12_0 m1_15755_n208# m1_16599_2028# m1_17703_788# vss nfet$12
Xnfet$14_3 m1_17926_34# vss m1_18496_1828# vss nfet$14
Xpfet$13_2 m1_n15602_4493# vdd vdd m1_n15602_4493# m1_n15874_4493# m1_n15874_4493#
+ m1_n15602_4493# vdd m1_n15874_4493# m1_n15874_4493# pfet$13
Xnfet$14_13 ref vss m1_16242_6960# vss nfet$14
Xpfet$7_6 m1_4402_7868# m1_4402_7868# m1_3254_4493# vdd m1_3254_4493# m1_4402_7868#
+ vdd vdd m1_3254_4493# m1_4402_7868# m1_3254_4493# m1_3254_4493# m1_4402_7868# m1_3254_4493#
+ vdd m1_3254_4493# vdd m1_3254_4493# pfet$7
Xpfet$5_3 vdd vdd m1_n1748_5099# m1_n2336_5099# pfet$5
Xpfet$9_11 vdd vdd m1_16599_5522# m1_15979_5220# pfet$9
Xnfet$6_0 m1_10834_1478# vss m1_11370_n340# vss nfet$6
Xnfet$14_4 m1_12790_n340# vss m1_15618_394# vss nfet$14
Xpfet$7_7 m1_8596_7868# m1_8596_7868# m1_7448_4493# vdd m1_7448_4493# m1_8596_7868#
+ vdd vdd m1_7448_4493# m1_8596_7868# m1_7448_4493# m1_7448_4493# m1_8596_7868# m1_7448_4493#
+ vdd m1_7448_4493# vdd m1_7448_4493# pfet$7
Xpfet$11_0 vdd m1_17926_34# vdd m1_17703_788# pfet$11
Xnfet$12_1 m1_15618_394# m1_16242_n208# m1_15979_2344# vss nfet$12
Xpfet$5_4 vdd vdd m1_6640_5099# m1_4402_7868# pfet$5
Xpfet$9_12 vdd vdd m1_16242_6960# ref pfet$9
Xnfet$6_1 m1_2446_1478# vss m1_2982_n340# vss nfet$6
Xnfet$12_2 m1_15618_394# m1_17703_788# m1_18496_1828# vss nfet$12
Xnfet$14_5 vss vss m1_17215_2028# vss nfet$14
Xpfet$11_1 vdd vdd m1_17926_34# m1_17215_2028# pfet$11
Xpfet$5_5 vdd vdd m1_10834_5099# m1_8596_7868# pfet$5
Xpfet$9_13 vdd vdd m1_15755_6960# m1_15618_7156# pfet$9
Xnfet$14_6 m1_17926_34# vss m1_19469_1832# vss nfet$14
Xnfet$6_2 m1_6640_1478# vss m1_7176_n340# vss nfet$6
Xpfet$11_2 vdd m1_16243_1828# vdd m1_17215_2028# pfet$11
Xnfet$12_3 m1_15755_n208# m1_15979_2344# m1_16243_1828# vss nfet$12
Xpfet$5_6 vdd vdd m1_2446_5099# m1_208_7868# pfet$5
Xnfet$10_0 m1_n7214_4493# vss m1_n7486_4493# m1_n7486_4493# m1_n7486_4493# m1_n7214_4493#
+ m1_n7214_4493# vss m1_n7486_4493# vss nfet$10
Xnfet$12_4 m1_15618_7156# m1_17703_6956# m1_18496_5840# vss nfet$12
Xnfet$6_3 m1_n1748_1478# vss m1_n1212_n340# vss nfet$6
Xnfet$14_7 vss vss m1_17215_5644# vss nfet$14
Xnfet$10_1 m1_n15602_4493# vss m1_n15874_4493# m1_n15874_4493# m1_n15874_4493# m1_n15602_4493#
+ m1_n15602_4493# vss m1_n15874_4493# vss nfet$10
Xpfet$11_3 vdd vdd m1_16243_1828# m1_16599_2028# pfet$11
Xpfet$5_7 vdd vdd m1_2446_1478# m1_208_n340# pfet$5
Xnfet$14_8 m1_17926_7472# vss m1_19469_4920# vss nfet$14
Xnfet$6_4 m1_10834_5099# vss m1_11370_4493# vss nfet$6
Xnfet$12_5 m1_15755_6960# m1_15979_5220# m1_16243_5840# vss nfet$12
Xnfet$10_2 m1_n11408_4493# vss m1_n11680_4493# m1_n11680_4493# m1_n11680_4493# m1_n11408_4493#
+ m1_n11408_4493# vss m1_n11680_4493# vss nfet$10
Xpfet$11_4 vdd m1_16243_5840# vdd m1_17215_5644# pfet$11
Xnfet$6_5 m1_6640_5099# vss m1_7176_4493# vss nfet$6
Xnfet$14_9 m1_17926_7472# vss m1_18496_5840# vss nfet$14
Xnfet$12_6 m1_15618_7156# m1_16242_6960# m1_15979_5220# vss nfet$12
Xpfet$11_5 vdd vdd m1_16243_5840# m1_16599_5522# pfet$11
Xnfet$6_6 m1_n1748_5099# vss m1_n1212_4493# vss nfet$6
Xnfet$12_7 m1_15755_6960# m1_16599_5522# m1_17703_6956# vss nfet$12
Xnfet$19_0 m1_19675_2344# vss lock vss nfet$19
Xpfet$11_6 vdd m1_17926_7472# vdd m1_17703_6956# pfet$11
Xnfet$6_7 m1_2446_5099# vss m1_2982_4493# vss nfet$6
Xpfet$11_7 vdd vdd m1_17926_7472# m1_17215_5644# pfet$11
Xpfet$18_0 vdd m1_19675_2344# vdd m1_19469_1832# pfet$18
Xpfet$18_1 vdd vdd m1_19675_2344# m1_19469_4920# pfet$18
.ends

.subckt nfet$31 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$32 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$31 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$32 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt xp_3_1_MUX S0 S1 VDD VSS OUT_1 C_1 B_1 A_1
Xnfet$31_2 S1 m1_239_n318# OUT_1 VSS nfet$31
Xnfet$31_3 S0 A_1 m1_239_n318# VSS nfet$31
Xnfet$32_0 S1 VSS m1_n432_n1290# VSS nfet$32
Xpfet$31_0 VDD A_1 m1_239_n318# m1_n432_458# pfet$31
Xnfet$32_1 S0 VSS m1_n432_458# VSS nfet$32
Xpfet$31_1 VDD C_1 OUT_1 S1 pfet$31
Xpfet$31_2 VDD B_1 m1_239_n318# S0 pfet$31
Xpfet$31_3 VDD m1_239_n318# OUT_1 m1_n432_n1290# pfet$31
Xpfet$32_0 VDD VDD m1_n432_n1290# S1 pfet$32
Xpfet$32_1 VDD VDD m1_n432_458# S0 pfet$32
Xnfet$31_1 m1_n432_458# B_1 m1_239_n318# VSS nfet$31
Xnfet$31_0 m1_n432_n1290# C_1 OUT_1 VSS nfet$31
.ends

.subckt nfet$20 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$25 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.5u
.ends

.subckt pfet$24 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$24 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt inv1u05u VDD in VSS out
Xpfet$24_0 VDD VDD out in pfet$24
Xnfet$24_0 in VSS out VSS nfet$24
.ends

.subckt pfet$22 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=4.55p ps=15.3u w=7u l=0.5u
.ends

.subckt nfet$22 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$21 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_954_0# w_n180_n88#
+ a_38_n60# a_n92_0# a_1058_n60# a_854_n60# a_342_0# a_138_0# a_650_n60#
X0 a_954_0# a_854_n60# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n60# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt pfet$23 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$23 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pass1u05u VDD VSS ind ins clkn clkp
Xpfet$23_0 VDD ind ins clkp pfet$23
Xnfet$23_0 clkn ind ins VSS nfet$23
.ends

.subckt nfet$21 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$20 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_954_0# w_n180_n88# a_854_n136#
+ a_n92_0# a_446_n136# a_650_n136# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt nfet$25 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt xp_programmable_basic_pump up vdd s1 s2 s3 s4 down out iref vss
Xnfet$20_10 pass1u05u_2/ins pass1u05u_2/ins m1_n7679_n8960# m1_n7679_n8960# out vss
+ nfet$20
Xpfet$25_3 vdd s4 pass1u05u_7/ins vdd pfet$25
Xinv1u05u_3 vdd s1 vss inv1u05u_3/out inv1u05u
Xnfet$20_11 vss vss vss vss vss vss nfet$20
Xpfet$22_20 vdd vdd vdd vdd pfet$22
Xnfet$20_12 down down vss vss m1_n7679_n8960# vss nfet$20
Xpfet$22_21 vdd vdd vdd vdd pfet$22
Xpfet$22_10 vdd vdd vdd vdd pfet$22
Xnfet$20_13 vss vss vss vss vss vss nfet$20
Xnfet$22_0 m1_n7879_n12170# pass1u05u_0/ins m1_n7879_n12170# out pass1u05u_0/ins vss
+ nfet$22
Xnfet$20_14 vss vss vss vss vss vss nfet$20
Xpfet$22_22 vdd vdd vdd vdd pfet$22
Xnfet$22_1 m1_n7879_n12170# pass1u05u_0/ins m1_n7879_n12170# out pass1u05u_0/ins vss
+ nfet$22
Xpfet$22_11 vdd vdd vdd vdd pfet$22
Xpfet$21_0 vdd vdd m1_n4127_3649# vss vss m1_n4127_3649# vdd vss vdd vss vss vdd m1_n4127_3649#
+ vss pfet$21
Xnfet$20_15 vss vss vss vss vss vss nfet$20
Xpfet$22_23 vdd vdd vdd vdd pfet$22
Xnfet$22_2 vss down vss m1_n7879_n12170# down vss nfet$22
Xpfet$21_1 m1_n5580_883# m1_n5580_883# out pass1u05u_5/ins pass1u05u_5/ins out vdd
+ pass1u05u_5/ins m1_n5580_883# pass1u05u_5/ins pass1u05u_5/ins m1_n5580_883# out
+ pass1u05u_5/ins pfet$21
Xpfet$22_12 vdd vdd vdd vdd pfet$22
Xpfet$22_13 vdd vdd vdd vdd pfet$22
Xnfet$22_3 vss down vss m1_n7879_n12170# down vss nfet$22
Xnfet$20_0 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out vss
+ nfet$20
Xpfet$21_2 m1_n5580_883# m1_n5580_883# out pass1u05u_5/ins pass1u05u_5/ins out vdd
+ pass1u05u_5/ins m1_n5580_883# pass1u05u_5/ins pass1u05u_5/ins m1_n5580_883# out
+ pass1u05u_5/ins pfet$21
Xpfet$22_14 vdd vdd vdd vdd pfet$22
Xnfet$22_4 vss down vss m1_n7879_n12170# down vss nfet$22
Xpfet$21_3 m1_n5580_883# m1_n5580_883# out pass1u05u_5/ins pass1u05u_5/ins out vdd
+ pass1u05u_5/ins m1_n5580_883# pass1u05u_5/ins pass1u05u_5/ins m1_n5580_883# out
+ pass1u05u_5/ins pfet$21
Xnfet$20_1 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out vss
+ nfet$20
Xpfet$22_15 vdd vdd vdd vdd pfet$22
Xnfet$22_5 vss down vss m1_n7879_n12170# down vss nfet$22
Xpfet$21_4 m1_n5580_883# m1_n5580_883# out pass1u05u_5/ins pass1u05u_5/ins out vdd
+ pass1u05u_5/ins m1_n5580_883# pass1u05u_5/ins pass1u05u_5/ins m1_n5580_883# out
+ pass1u05u_5/ins pfet$21
Xnfet$20_2 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out vss
+ nfet$20
Xpfet$22_16 vdd vdd vdd vdd pfet$22
Xnfet$22_6 m1_n7879_n12170# pass1u05u_0/ins m1_n7879_n12170# out pass1u05u_0/ins vss
+ nfet$22
Xpfet$21_5 m1_n4127_3649# m1_n4127_3649# pass1u05u_7/ind pass1u05u_7/ind pass1u05u_7/ind
+ pass1u05u_7/ind vdd pass1u05u_7/ind m1_n4127_3649# pass1u05u_7/ind pass1u05u_7/ind
+ m1_n4127_3649# pass1u05u_7/ind pass1u05u_7/ind pfet$21
Xnfet$20_3 vss vss vss vss vss vss nfet$20
Xpfet$22_17 vdd vdd vdd vdd pfet$22
Xnfet$20_4 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out vss
+ nfet$20
Xnfet$22_7 m1_n7879_n12170# pass1u05u_0/ins m1_n7879_n12170# out pass1u05u_0/ins vss
+ nfet$22
Xpfet$22_18 vdd vdd vdd vdd pfet$22
Xpass1u05u_0 vdd vss iref pass1u05u_0/ins s3 inv1u05u_1/out pass1u05u
Xnfet$22_8 vss vdd vss m1_n8144_n9165# vdd vss nfet$22
Xnfet$20_5 vss vss vss vss vss vss nfet$20
Xpfet$22_19 vdd vdd vdd vdd pfet$22
Xpass1u05u_1 vdd vss iref pass1u05u_1/ins s2 inv1u05u_2/out pass1u05u
Xnfet$20_6 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out vss
+ nfet$20
Xnfet$22_9 m1_n7216_n8262# iref m1_n7216_n8262# pass1u05u_7/ind iref vss nfet$22
Xnfet$21_10 vss vss vss vss vss vss nfet$21
Xpass1u05u_2 vdd vss iref pass1u05u_2/ins s1 inv1u05u_3/out pass1u05u
Xnfet$21_11 vss vss vss vss vss vss nfet$21
Xnfet$20_7 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out vss
+ nfet$20
Xpfet$20_20 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$20
Xpass1u05u_3 vdd vss pass1u05u_7/ind pass1u05u_3/ins s1 inv1u05u_3/out pass1u05u
Xnfet$20_8 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out vss
+ nfet$20
Xnfet$21_12 vss vss vss vss vss vss nfet$21
Xpfet$20_21 m1_n6703_2564# m1_n6703_2564# pass1u05u_4/ins out out vdd pass1u05u_4/ins
+ m1_n6703_2564# pass1u05u_4/ins pass1u05u_4/ins m1_n6703_2564# out pass1u05u_4/ins
+ pass1u05u_4/ins pfet$20
Xpfet$20_10 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$20
Xpass1u05u_4 vdd vss pass1u05u_7/ind pass1u05u_4/ins s2 inv1u05u_2/out pass1u05u
Xnfet$20_9 pass1u05u_6/ins pass1u05u_6/ins m1_n8807_n11192# m1_n8807_n11192# out vss
+ nfet$20
Xnfet$21_13 vss vss vss vss vss vss nfet$21
Xpfet$20_22 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$20
Xpfet$20_11 vdd vdd up m1_n5450_4559# m1_n5450_4559# vdd up vdd up up vdd m1_n5450_4559#
+ up up pfet$20
Xpass1u05u_5 vdd vss pass1u05u_7/ind pass1u05u_5/ins s3 inv1u05u_1/out pass1u05u
Xnfet$25_0 inv1u05u_2/out pass1u05u_1/ins vss vss nfet$25
Xpfet$20_23 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$20
Xpfet$20_12 vdd vdd up m1_n6703_2564# m1_n6703_2564# vdd up vdd up up vdd m1_n6703_2564#
+ up up pfet$20
Xpass1u05u_6 vdd vss iref pass1u05u_6/ins s4 inv1u05u_0/out pass1u05u
Xnfet$25_1 inv1u05u_3/out pass1u05u_2/ins vss vss nfet$25
Xpfet$20_24 m1_n5450_4559# m1_n5450_4559# pass1u05u_3/ins out out vdd pass1u05u_3/ins
+ m1_n5450_4559# pass1u05u_3/ins pass1u05u_3/ins m1_n5450_4559# out pass1u05u_3/ins
+ pass1u05u_3/ins pfet$20
Xpfet$20_13 vdd vdd up m1_n6703_2564# m1_n6703_2564# vdd up vdd up up vdd m1_n6703_2564#
+ up up pfet$20
Xpass1u05u_7 vdd vss pass1u05u_7/ind pass1u05u_7/ins s4 inv1u05u_0/out pass1u05u
Xnfet$25_2 inv1u05u_0/out pass1u05u_6/ins vss vss nfet$25
Xpfet$20_25 m1_n6703_2564# m1_n6703_2564# pass1u05u_4/ins out out vdd pass1u05u_4/ins
+ m1_n6703_2564# pass1u05u_4/ins pass1u05u_4/ins m1_n6703_2564# out pass1u05u_4/ins
+ pass1u05u_4/ins pfet$20
Xpfet$20_14 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$20
Xnfet$25_3 inv1u05u_1/out pass1u05u_0/ins vss vss nfet$25
Xpfet$20_15 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$20
Xpfet$22_0 vdd vdd vdd vdd pfet$22
Xpfet$20_16 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$20
Xpfet$20_17 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$20
Xpfet$22_1 vdd vdd vdd vdd pfet$22
Xpfet$20_18 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$20
Xnfet$21_0 down down vss vss m1_n8807_n11192# vss nfet$21
Xpfet$22_2 vdd vdd vdd vdd pfet$22
Xpfet$20_19 m1_n8156_628# m1_n8156_628# pass1u05u_7/ins out out vdd pass1u05u_7/ins
+ m1_n8156_628# pass1u05u_7/ins pass1u05u_7/ins m1_n8156_628# out pass1u05u_7/ins
+ pass1u05u_7/ins pfet$20
Xnfet$21_1 down down vss vss m1_n8807_n11192# vss nfet$21
Xpfet$22_3 vdd vdd vdd vdd pfet$22
Xpfet$20_0 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$20
Xnfet$21_2 down down vss vss m1_n8807_n11192# vss nfet$21
Xnfet$22_10 m1_n8607_n8040# pass1u05u_1/ins m1_n8607_n8040# out pass1u05u_1/ins vss
+ nfet$22
Xpfet$22_4 vdd vdd vdd vdd pfet$22
Xpfet$20_1 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$20
Xnfet$21_3 down down vss vss m1_n8807_n11192# vss nfet$21
Xnfet$22_11 m1_n8144_n9165# iref m1_n8144_n9165# iref iref vss nfet$22
Xpfet$22_5 vdd vdd vdd vdd pfet$22
Xpfet$20_2 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$20
Xnfet$22_12 vss down vss m1_n8607_n8040# down vss nfet$22
Xpfet$22_6 vdd vdd vdd vdd pfet$22
Xnfet$21_4 vss vss vss vss vss vss nfet$21
Xpfet$20_3 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$20
Xnfet$21_5 vss vss vss vss vss vss nfet$21
Xnfet$22_13 vss vdd vss m1_n7216_n8262# vdd vss nfet$22
Xpfet$22_7 vdd vdd vdd vdd pfet$22
Xpfet$20_4 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$20
Xnfet$22_14 m1_n8607_n8040# pass1u05u_1/ins m1_n8607_n8040# out pass1u05u_1/ins vss
+ nfet$22
Xnfet$21_6 down down vss vss m1_n8807_n11192# vss nfet$21
Xpfet$20_5 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$20
Xpfet$22_8 vdd vdd vdd vdd pfet$22
Xnfet$21_7 down down vss vss m1_n8807_n11192# vss nfet$21
Xnfet$22_15 vss down vss m1_n8607_n8040# down vss nfet$22
Xpfet$22_9 vdd vdd vdd vdd pfet$22
Xpfet$20_6 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$20
Xnfet$21_8 down down vss vss m1_n8807_n11192# vss nfet$21
Xpfet$20_7 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$20
Xnfet$21_9 down down vss vss m1_n8807_n11192# vss nfet$21
Xpfet$20_8 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$20
Xpfet$20_9 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$20
Xpfet$25_0 vdd s3 pass1u05u_5/ins vdd pfet$25
Xinv1u05u_0 vdd s4 vss inv1u05u_0/out inv1u05u
Xpfet$25_1 vdd s2 pass1u05u_4/ins vdd pfet$25
Xinv1u05u_1 vdd s3 vss inv1u05u_1/out inv1u05u
Xpfet$25_2 vdd s1 pass1u05u_3/ins vdd pfet$25
Xinv1u05u_2 vdd s2 vss inv1u05u_2/out inv1u05u
.ends

.subckt nfet$55 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$54 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt asc_delay vdd in vss out
Xnfet$55_0 m1_878_n53# vss out vss nfet$55
Xnfet$55_1 in vss m1_878_n53# vss nfet$55
Xpfet$54_0 vdd vdd out m1_878_n53# pfet$54
Xpfet$54_1 vdd vdd m1_878_n53# in pfet$54
.ends

.subckt pfet$39 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$45 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt nfet$38 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt pfet$44 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt pfet$37 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$43 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$42 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$36 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$35 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$41 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt nfet$34 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$40 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$33 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$46 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$45 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$39 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$38 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt nfet$44 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt pfet$43 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt nfet$37 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$36 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$42 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$35 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$41 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt pfet$34 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$40 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$33 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_PFD_DFF_20250831 vss fref down up vdd fdiv
Xpfet$39_0 vdd vdd m1_n3885_n4045# m1_n5428_n3533# pfet$39
Xnfet$45_0 m1_n4677_n8889# m1_n1925_n10720# vss vss nfet$45
Xpfet$39_1 vdd vdd m1_n5650_n4045# m1_n5868_n3849# pfet$39
Xnfet$45_1 m1_n1925_n10720# m1_n3098_n10720# vss vss nfet$45
Xnfet$38_0 m1_n1926_n4095# m1_n3099_n4095# vss vss nfet$38
Xpfet$39_2 vdd vdd m1_n3885_n6084# m1_n5428_n5842# pfet$39
Xpfet$44_0 m1_n4677_n8889# vdd vdd m1_n1925_n10720# pfet$44
Xpfet$44_1 m1_n1925_n10720# vdd vdd m1_n3098_n10720# pfet$44
Xnfet$45_2 m1_n4677_n10522# m1_n1925_n9135# vss vss nfet$45
Xnfet$38_1 m1_n4678_n3849# m1_n1926_n5680# vss vss nfet$38
Xpfet$39_3 vdd vdd m1_n5868_n3849# fref pfet$39
Xpfet$37_0 vdd vdd m1_5464_n5483# m1_5895_n8089# pfet$37
Xnfet$45_3 m1_n1925_n9135# m1_n3098_n9135# vss vss nfet$45
Xnfet$38_2 m1_n1926_n5680# m1_n3099_n5680# vss vss nfet$38
Xnfet$43_0 m1_n3884_n9085# m1_1095_n11125# m1_832_n8573# vss nfet$43
Xpfet$44_2 m1_n4677_n10522# vdd vdd m1_n1925_n9135# pfet$44
Xpfet$37_1 vdd vdd m1_4978_n5483# m1_5464_n5483# pfet$37
Xpfet$44_3 m1_n1925_n9135# vdd vdd m1_n3098_n9135# pfet$44
Xnfet$38_3 m1_n4678_n5482# m1_n1926_n4095# vss vss nfet$38
Xpfet$42_0 vdd vdd m1_2779_n10883# m1_2068_n8889# pfet$42
Xnfet$43_1 m1_n3884_n11124# m1_1452_n8889# m1_2556_n10129# vss nfet$43
Xnfet$36_0 m1_4978_n5483# vss m1_2758_n8889# vss nfet$36
Xnfet$43_2 m1_832_n8573# vss m1_1452_n8889# vss nfet$43
Xpfet$42_1 vdd m1_2779_n10883# vdd m1_2556_n10129# pfet$42
Xpfet$35_0 vdd vdd m1_3349_n5165# m1_2779_n3533# pfet$35
Xpfet$42_2 vdd m1_1095_n11125# m1_832_n8573# m1_n3884_n11124# pfet$42
Xnfet$43_3 vdd vss m1_1095_n11125# vss nfet$43
Xnfet$41_0 m1_n3885_n4045# vss m1_n3099_n4095# vss nfet$41
Xpfet$35_1 vdd vdd up m1_2779_n3533# pfet$35
Xnfet$43_4 m1_n3884_n11124# m1_832_n8573# m1_1096_n9089# vss nfet$43
Xnfet$34_0 m1_2068_n5361# m1_2068_n5361# vss vss m1_1550_n5165# vss nfet$34
Xpfet$35_2 vdd vdd m1_2068_n5361# m1_2758_n8889# pfet$35
Xpfet$42_3 vdd m1_1452_n8889# m1_2556_n10129# m1_n3884_n9085# pfet$42
Xnfet$41_1 m1_n3885_n6084# vss m1_n3099_n5680# vss nfet$41
Xpfet$40_0 vdd m1_n5428_n3533# vdd m1_n5650_n4045# pfet$40
Xpfet$35_3 vdd vdd m1_1452_n5483# m1_832_n5785# pfet$35
Xnfet$34_1 m1_1452_n5483# m1_1452_n5483# m1_1096_n5165# m1_1096_n5165# m1_1550_n5165#
+ vss nfet$34
Xpfet$42_4 vdd vdd m1_1452_n8889# m1_832_n8573# pfet$42
Xnfet$43_5 m1_2758_n8889# vss m1_2068_n8889# vss nfet$43
Xpfet$33_0 vdd m1_832_n5785# m1_1096_n5165# m1_n3885_n6084# pfet$33
Xpfet$40_1 vdd vdd m1_n5428_n3533# m1_n4678_n3849# pfet$40
Xnfet$43_6 m1_2779_n10883# vss down vss nfet$43
Xpfet$35_4 vdd vdd m1_1095_n4045# vdd pfet$35
Xnfet$34_2 m1_2556_n4049# m1_2556_n4049# vss vss m1_3015_n4205# vss nfet$34
Xpfet$42_5 vdd vdd m1_1095_n11125# vdd pfet$42
Xpfet$33_1 vdd m1_1452_n5483# m1_2556_n4049# m1_n3885_n6084# pfet$33
Xpfet$40_2 vdd m1_n5428_n5842# vdd m1_n5868_n3849# pfet$40
Xnfet$43_10 m1_n5867_n10544# vss m1_n5649_n11124# vss nfet$43
Xnfet$34_3 m1_2068_n5361# m1_2068_n5361# m1_2779_n3533# m1_2779_n3533# m1_3015_n4205#
+ vss nfet$34
Xpfet$42_6 vdd vdd m1_1096_n9089# m1_1452_n8889# pfet$42
Xnfet$43_7 m1_2779_n10883# vss m1_3349_n9089# vss nfet$43
Xpfet$33_2 vdd m1_1095_n4045# m1_832_n5785# m1_n3885_n4045# pfet$33
Xpfet$40_3 vdd vdd m1_n5428_n5842# m1_n4678_n5482# pfet$40
Xnfet$43_11 fdiv vss m1_n5867_n10544# vss nfet$43
Xnfet$43_8 m1_n3884_n9085# m1_2556_n10129# m1_3349_n9089# vss nfet$43
Xpfet$42_20 vdd m1_n5427_n8573# vdd m1_n5867_n10544# pfet$42
Xpfet$42_7 vdd m1_832_n8573# m1_1096_n9089# m1_n3884_n9085# pfet$42
Xpfet$33_3 vdd m1_2556_n4049# m1_3349_n5165# m1_n3885_n4045# pfet$33
Xnfet$43_12 m1_n5427_n8573# vss m1_n3884_n9085# vss nfet$43
Xpfet$42_10 vdd vdd m1_3349_n9089# m1_2779_n10883# pfet$42
Xnfet$43_9 m1_n5427_n10882# vss m1_n3884_n11124# vss nfet$43
Xpfet$42_8 vdd m1_1096_n9089# vdd m1_2068_n8889# pfet$42
Xpfet$42_11 vdd vdd down m1_2779_n10883# pfet$42
Xpfet$42_9 vdd vdd m1_2068_n8889# m1_2758_n8889# pfet$42
Xpfet$42_12 vdd m1_2556_n10129# m1_3349_n9089# m1_n3884_n11124# pfet$42
Xpfet$42_13 vdd vdd m1_n5427_n8573# m1_n4677_n8889# pfet$42
Xpfet$42_14 vdd vdd m1_n3884_n11124# m1_n5427_n10882# pfet$42
Xnfet$46_0 up up m1_5895_n8089# m1_5895_n8089# m1_5043_n9245# vss nfet$46
Xpfet$42_15 vdd m1_n5427_n10882# vdd m1_n5649_n11124# pfet$42
Xpfet$45_0 vdd m1_5895_n8089# vdd down pfet$45
Xnfet$46_1 down down vss vss m1_5043_n9245# vss nfet$46
Xnfet$39_0 m1_n5428_n3533# vss m1_n3885_n4045# vss nfet$39
Xpfet$42_16 vdd vdd m1_n5427_n10882# m1_n4677_n10522# pfet$42
Xnfet$39_1 m1_n5868_n3849# vss m1_n5650_n4045# vss nfet$39
Xpfet$45_1 vdd vdd m1_5895_n8089# up pfet$45
Xpfet$38_0 m1_n1926_n4095# vdd vdd m1_n3099_n4095# pfet$38
Xpfet$42_17 vdd vdd m1_n5649_n11124# m1_n5867_n10544# pfet$42
Xnfet$44_0 m1_n3884_n11124# vss m1_n3098_n10720# vss nfet$44
Xpfet$38_1 m1_n4678_n3849# vdd vdd m1_n1926_n5680# pfet$38
Xnfet$39_2 m1_n5428_n5842# vss m1_n3885_n6084# vss nfet$39
Xpfet$42_18 vdd vdd m1_n5867_n10544# fdiv pfet$42
Xnfet$39_3 fref vss m1_n5868_n3849# vss nfet$39
Xpfet$43_0 vdd vdd m1_n3098_n10720# m1_n3884_n11124# pfet$43
Xnfet$44_1 m1_n3884_n9085# vss m1_n3098_n9135# vss nfet$44
Xpfet$38_2 m1_n1926_n5680# vdd vdd m1_n3099_n5680# pfet$38
Xnfet$37_0 m1_5895_n8089# vss m1_5464_n5483# vss nfet$37
Xpfet$42_19 vdd vdd m1_n3884_n9085# m1_n5427_n8573# pfet$42
Xpfet$38_3 m1_n4678_n5482# vdd vdd m1_n1926_n4095# pfet$38
Xnfet$37_1 m1_5464_n5483# vss m1_4978_n5483# vss nfet$37
Xpfet$43_1 vdd vdd m1_n3098_n9135# m1_n3884_n9085# pfet$43
Xpfet$36_0 vdd vdd m1_2758_n8889# m1_4978_n5483# pfet$36
Xnfet$42_0 m1_2556_n10129# m1_2556_n10129# vss vss m1_3015_n10205# vss nfet$42
Xnfet$42_1 m1_1452_n8889# m1_1452_n8889# m1_1096_n9089# m1_1096_n9089# m1_1550_n9245#
+ vss nfet$42
Xnfet$35_0 m1_2779_n3533# vss up vss nfet$35
Xpfet$41_0 vdd vdd m1_n3099_n4095# m1_n3885_n4045# pfet$41
Xpfet$34_0 vdd vdd m1_1096_n5165# m1_1452_n5483# pfet$34
Xnfet$42_2 m1_2068_n8889# m1_2068_n8889# vss vss m1_1550_n9245# vss nfet$42
Xpfet$41_1 vdd vdd m1_n3099_n5680# m1_n3885_n6084# pfet$41
Xnfet$35_1 m1_2779_n3533# vss m1_3349_n5165# vss nfet$35
Xnfet$35_2 m1_2758_n8889# vss m1_2068_n5361# vss nfet$35
Xnfet$42_3 m1_2068_n8889# m1_2068_n8889# m1_2779_n10883# m1_2779_n10883# m1_3015_n10205#
+ vss nfet$42
Xpfet$34_1 vdd m1_1096_n5165# vdd m1_2068_n5361# pfet$34
Xnfet$40_0 m1_n4678_n3849# m1_n4678_n3849# m1_n5428_n3533# m1_n5428_n3533# m1_n5192_n4205#
+ vss nfet$40
Xnfet$35_3 m1_832_n5785# vss m1_1452_n5483# vss nfet$35
Xpfet$34_2 vdd m1_2779_n3533# vdd m1_2556_n4049# pfet$34
Xnfet$42_4 m1_n4677_n10522# m1_n4677_n10522# m1_n5427_n10882# m1_n5427_n10882# m1_n5191_n10204#
+ vss nfet$42
Xnfet$40_1 m1_n5650_n4045# m1_n5650_n4045# vss vss m1_n5192_n4205# vss nfet$40
Xnfet$33_0 m1_n3885_n4045# m1_832_n5785# m1_1096_n5165# vss nfet$33
Xnfet$35_4 vdd vss m1_1095_n4045# vss nfet$35
Xnfet$42_5 m1_n5649_n11124# m1_n5649_n11124# vss vss m1_n5191_n10204# vss nfet$42
Xpfet$34_3 vdd vdd m1_2779_n3533# m1_2068_n5361# pfet$34
Xnfet$33_1 m1_n3885_n4045# m1_1452_n5483# m1_2556_n4049# vss nfet$33
Xnfet$40_2 m1_n4678_n5482# m1_n4678_n5482# m1_n5428_n5842# m1_n5428_n5842# m1_n5192_n5164#
+ vss nfet$40
Xnfet$42_6 m1_n4677_n8889# m1_n4677_n8889# m1_n5427_n8573# m1_n5427_n8573# m1_n5191_n9245#
+ vss nfet$42
Xnfet$33_2 m1_n3885_n6084# m1_1095_n4045# m1_832_n5785# vss nfet$33
Xnfet$40_3 m1_n5868_n3849# m1_n5868_n3849# vss vss m1_n5192_n5164# vss nfet$40
Xnfet$42_7 m1_n5867_n10544# m1_n5867_n10544# vss vss m1_n5191_n9245# vss nfet$42
Xnfet$33_3 m1_n3885_n6084# m1_2556_n4049# m1_3349_n5165# vss nfet$33
.ends

.subckt nfet$54 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$53 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$52 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.5u
.ends

.subckt pfet$51 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=9.75p pd=31.3u as=9.75p ps=31.3u w=15u l=0.5u
.ends

.subckt cap_mim m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
.ends

.subckt nfet$53 a_n84_0# a_38_n132# a_138_0# VSUBS
X0 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.5u
.ends

.subckt pfet$52 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=9.75p pd=31.3u as=9.75p ps=31.3u w=15u l=0.5u
.ends

.subckt CSRVCO_20250823 vctrl vosc vdd vss
Xnfet$54_0 m1_n8380_274# vss vosc vss nfet$54
Xpfet$53_0 vdd vdd vosc m1_n8380_274# pfet$53
Xnfet$54_1 m1_n11916_1270# vss m1_n8380_274# vss nfet$54
Xpfet$53_1 vdd vdd m1_n8380_274# m1_n11916_1270# pfet$53
Xnfet$52_0 m1_n9838_266# m1_n12754_674# m1_n9352_266# vss nfet$52
Xpfet$51_0 vdd vdd m1_n12264_2422# m1_n16019_266# pfet$51
Xnfet$52_1 vctrl vss m1_n12268_985# vss nfet$52
Xpfet$51_1 vdd vdd m1_n14208_3657# m1_n16019_266# pfet$51
Xnfet$52_2 vctrl vss m1_n14283_186# vss nfet$52
Xpfet$51_2 vdd vdd m1_n13722_3340# m1_n16019_266# pfet$51
Xnfet$52_3 vctrl vss m1_n13794_186# vss nfet$52
Xnfet$52_4 vctrl vss m1_n13240_368# vss nfet$52
Xpfet$51_4 vdd vdd m1_n13236_3035# m1_n16019_266# pfet$51
Xpfet$51_3 vdd m1_n16019_266# vdd m1_n16019_266# pfet$51
Xnfet$52_5 vctrl vss m1_n12754_674# vss nfet$52
Xpfet$51_5 vdd vdd m1_n14693_3963# m1_n16019_266# pfet$51
Xcap_mim_0 vss m1_n11296_266# cap_mim
Xnfet$52_6 vctrl m1_n16019_266# vss vss nfet$52
Xpfet$51_6 vdd vdd m1_n12750_2729# m1_n16019_266# pfet$51
Xcap_mim_1 vss m1_n10810_266# cap_mim
Xnfet$52_7 vctrl vss m1_n15245_186# vss nfet$52
Xpfet$51_7 vdd vdd m1_n15180_4275# m1_n16019_266# pfet$51
Xcap_mim_2 vss m1_n10324_266# cap_mim
Xnfet$52_8 vctrl vss m1_n14765_186# vss nfet$52
Xpfet$51_8 vdd m1_n13236_3035# m1_n9838_266# m1_n10324_266# pfet$51
Xnfet$52_9 m1_n10324_266# m1_n13240_368# m1_n9838_266# vss nfet$52
Xcap_mim_3 vss m1_n11916_1270# cap_mim
Xpfet$51_9 vdd m1_n12750_2729# m1_n9352_266# m1_n9838_266# pfet$51
Xcap_mim_5 vss m1_n9838_266# cap_mim
Xcap_mim_4 vss m1_n9352_266# cap_mim
Xcap_mim_6 vss m1_n11782_266# cap_mim
Xnfet$53_0 vss vss vss vss nfet$53
Xnfet$53_1 vss vss vss vss nfet$53
Xpfet$52_1 vdd vdd vdd vdd pfet$52
Xpfet$52_0 vdd vdd vdd vdd pfet$52
Xnfet$52_10 m1_n9352_266# m1_n12268_985# m1_n11916_1270# vss nfet$52
Xnfet$52_11 m1_n11916_1270# m1_n15245_186# m1_n11782_266# vss nfet$52
Xpfet$51_10 vdd m1_n14208_3657# m1_n10810_266# m1_n11296_266# pfet$51
Xnfet$52_12 m1_n11782_266# m1_n14765_186# m1_n11296_266# vss nfet$52
Xpfet$51_11 vdd m1_n12264_2422# m1_n11916_1270# m1_n9352_266# pfet$51
Xnfet$52_13 m1_n11296_266# m1_n14283_186# m1_n10810_266# vss nfet$52
Xnfet$52_14 m1_n10810_266# m1_n13794_186# m1_n10324_266# vss nfet$52
Xpfet$51_12 vdd m1_n14693_3963# m1_n11296_266# m1_n11782_266# pfet$51
Xpfet$51_13 vdd m1_n13722_3340# m1_n10324_266# m1_n10810_266# pfet$51
Xpfet$51_14 vdd m1_n15180_4275# m1_n11782_266# m1_n11916_1270# pfet$51
.ends

.subckt top_level_nosc_20250831 div_def div_prc_s8 div_prc_s7 div_prc_s6 div_prc_s5
+ div_prc_s4 div_prc_s3 div_prc_s2 div_prc_s1 div_prc_s0 div_out div_in div_swc_s0
+ div_swc_s1 div_swc_s2 div_swc_s3 div_swc_s4 div_swc_s5 div_swc_s6 div_swc_s7 div_swc_s8
+ lock ref ext_pfd_div ext_pfd_ref ext_pfd_up ext_pfd_down mx_pfd_s1 mx_pfd_s0 up
+ down cp_s1 cp_s2 cp_s3 cp_s4 i_cp_100u filter_in out filter_out ext_vco_in ext_vco_out
+ mx_vco_s0 mx_vco_s1 vdd vss
Xasc_drive_buffer_up_0 vss vdd asc_drive_buffer_up_0/out xp_3_1_MUX_5/OUT_1 asc_drive_buffer_up
Xasc_dual_psd_def_20250809_0 asc_dual_psd_def_20250809_0/vdd vss div_prc_s0 div_prc_s1
+ div_prc_s2 div_prc_s3 div_prc_s4 div_prc_s5 div_prc_s6 div_prc_s7 div_prc_s8 xp_3_1_MUX_3/OUT_1
+ div_swc_s0 div_swc_s1 div_swc_s2 div_swc_s3 div_swc_s4 div_swc_s5 div_swc_s6 div_swc_s7
+ div_swc_s8 asc_delay_0/out div_def vdd asc_dual_psd_def_20250809
Xasc_drive_buffer_0 vss asc_delay_0/in vdd out asc_drive_buffer
Xasc_drive_buffer_1 vss asc_delay_0/out vdd div_in asc_drive_buffer
Xasc_drive_buffer_2 vss xp_3_1_MUX_3/OUT_1 vdd div_out asc_drive_buffer
Xasc_drive_buffer_3 vss xp_3_1_MUX_5/OUT_1 vdd up asc_drive_buffer
Xasc_hysteresis_buffer_0 vss ref vdd xp_3_1_MUX_2/OUT_1 asc_hysteresis_buffer
Xasc_drive_buffer_4 vss xp_3_1_MUX_4/OUT_1 vdd down asc_drive_buffer
Xasc_lock_detector_20250826_0 xp_3_1_MUX_2/OUT_1 vdd xp_3_1_MUX_3/OUT_1 asc_drive_buffer_6/in
+ vss asc_lock_detector_20250826
Xasc_drive_buffer_5 vss xp_3_1_MUX_4/OUT_1 vdd asc_drive_buffer_5/out asc_drive_buffer
Xasc_drive_buffer_6 vss asc_drive_buffer_6/in vdd lock asc_drive_buffer
Xxp_3_1_MUX_0 mx_vco_s0 mx_vco_s1 vdd vss asc_delay_0/in xp_3_1_MUX_0/C_1 xp_3_1_MUX_0/B_1
+ ext_vco_out xp_3_1_MUX
Xxp_3_1_MUX_1 mx_vco_s0 mx_vco_s1 vdd vss filter_out xp_3_1_MUX_1/C_1 xp_3_1_MUX_1/B_1
+ ext_vco_in xp_3_1_MUX
Xxp_3_1_MUX_2 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX_2/OUT_1 xp_3_1_MUX_2/C_1 xp_3_1_MUX_2/B_1
+ ext_pfd_ref xp_3_1_MUX
Xxp_3_1_MUX_3 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX_3/OUT_1 xp_3_1_MUX_3/C_1 xp_3_1_MUX_3/B_1
+ ext_pfd_div xp_3_1_MUX
Xxp_3_1_MUX_4 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX_4/OUT_1 xp_3_1_MUX_4/C_1 xp_3_1_MUX_4/B_1
+ ext_pfd_down xp_3_1_MUX
Xxp_3_1_MUX_5 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX_5/OUT_1 xp_3_1_MUX_5/C_1 xp_3_1_MUX_5/B_1
+ ext_pfd_up xp_3_1_MUX
Xxp_programmable_basic_pump_0 asc_drive_buffer_up_0/out vdd cp_s1 cp_s2 cp_s3 cp_s4
+ asc_drive_buffer_5/out filter_in i_cp_100u vss xp_programmable_basic_pump
Xasc_delay_0 vdd asc_delay_0/in vss asc_delay_0/out asc_delay
Xasc_PFD_DFF_20250831_0 vss xp_3_1_MUX_2/C_1 xp_3_1_MUX_4/C_1 xp_3_1_MUX_5/C_1 vdd
+ xp_3_1_MUX_3/C_1 asc_PFD_DFF_20250831
Xasc_PFD_DFF_20250831_1 vss xp_3_1_MUX_2/B_1 xp_3_1_MUX_5/B_1 xp_3_1_MUX_4/B_1 vdd
+ xp_3_1_MUX_3/B_1 asc_PFD_DFF_20250831
XCSRVCO_20250823_0 xp_3_1_MUX_1/C_1 xp_3_1_MUX_0/C_1 vdd vss CSRVCO_20250823
.ends

