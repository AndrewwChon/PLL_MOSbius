* Extracted by KLayout with GF180MCU LVS runset on : 29/07/2025 04:22

.SUBCKT pass1u05u vss clkn ind ins vdd clkp
M$1 ins clkp ind vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$2 ins clkn ind vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
.ENDS pass1u05u
