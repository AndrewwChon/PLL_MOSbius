* NGSPICE file created from VCOfinal_noCP.ext - technology: gf180mcuD

.subckt nfet$19$1 a_30_260# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_260# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$6 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=1.625p ps=6.3u w=2.5u l=0.28u
.ends

.subckt pfet$4 a_1054_0# a_734_0# a_254_0# a_894_0# a_348_560# a_828_560# a_988_560#
+ w_n180_n88# a_1214_0# a_414_0# a_n92_0# a_94_0# a_574_0# a_508_560# a_188_560# a_668_560#
+ a_1148_560# a_28_560#
X0 a_1214_0# a_1148_560# a_1054_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_734_0# a_668_560# a_574_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X3 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X4 a_1054_0# a_988_560# a_894_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X5 a_894_0# a_828_560# a_734_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X6 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X7 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$5 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt pfet$5 a_254_0# a_348_560# w_n180_n88# a_414_0# a_n92_0# a_94_0# a_574_0#
+ a_508_560# a_188_560# a_28_560#
X0 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$6 a_254_0# a_n84_0# a_94_0# a_190_460# a_30_460# VSUBS
X0 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt nfet$4 a_1054_0# a_734_0# a_510_n132# a_254_0# a_894_0# a_670_n132# a_1214_0#
+ a_830_n132# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132# a_574_0# a_990_n132#
+ a_350_n132# a_1150_n132# VSUBS
X0 a_734_0# a_670_n132# a_574_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X3 a_1054_0# a_990_n132# a_894_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X4 a_894_0# a_830_n132# a_734_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X5 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X6 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X7 a_1214_0# a_1150_n132# a_1054_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt Pcomparator vss vdd iref inn inp out
Xpfet$6_0 vdd vdd vdd vdd pfet$6
Xpfet$6_2 vdd vdd vdd vdd pfet$6
Xpfet$6_1 vdd vdd vdd vdd pfet$6
Xpfet$4_0 out out vdd vdd iref iref iref vdd vdd out vdd out vdd iref iref iref iref
+ iref pfet$4
Xpfet$6_3 vdd vdd vdd vdd pfet$6
Xpfet$4_1 out out vdd vdd iref iref iref vdd vdd out vdd out vdd iref iref iref iref
+ iref pfet$4
Xnfet$5_0 vss vss vss vss vss vss vss vss vss vss nfet$5
Xnfet$5_1 vss vss vss vss vss vss vss vss vss vss nfet$5
Xpfet$5_10 vdd iref vdd iref vdd iref vdd iref iref iref pfet$5
Xpfet$5_12 m1_2779_n1752# inn vdd m1_3615_n1223# m1_2779_n1752# m1_3615_n1223# m1_2779_n1752#
+ inn inn inn pfet$5
Xpfet$5_11 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$5
Xpfet$5_13 m1_2779_n1752# inp vdd m1_5539_n2811# m1_2779_n1752# m1_5539_n2811# m1_2779_n1752#
+ inp inp inp pfet$5
Xpfet$5_0 m1_2779_n1752# inp vdd m1_5539_n2811# m1_2779_n1752# m1_5539_n2811# m1_2779_n1752#
+ inp inp inp pfet$5
Xpfet$5_1 m1_2779_n1752# m1_2779_n1752# vdd m1_2779_n1752# m1_2779_n1752# m1_2779_n1752#
+ m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# pfet$5
Xpfet$5_2 m1_2779_n1752# inn vdd m1_3615_n1223# m1_2779_n1752# m1_3615_n1223# m1_2779_n1752#
+ inn inn inn pfet$5
Xpfet$5_3 m1_2779_n1752# m1_2779_n1752# vdd m1_2779_n1752# m1_2779_n1752# m1_2779_n1752#
+ m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# pfet$5
Xnfet$6_0 vss vss m1_3615_n1223# m1_3615_n1223# m1_3615_n1223# vss nfet$6
Xpfet$5_4 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$5
Xnfet$6_1 vss vss m1_5539_n2811# m1_3615_n1223# m1_3615_n1223# vss nfet$6
Xpfet$5_6 vdd iref vdd iref vdd iref vdd iref iref iref pfet$5
Xpfet$5_5 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$5
Xnfet$6_2 vss vss m1_5539_n2811# m1_3615_n1223# m1_3615_n1223# vss nfet$6
Xnfet$4_0 out out m1_5539_n2811# vss vss m1_5539_n2811# vss m1_5539_n2811# out m1_5539_n2811#
+ vss out m1_5539_n2811# vss m1_5539_n2811# m1_5539_n2811# m1_5539_n2811# vss nfet$4
Xpfet$5_7 vdd iref vdd iref vdd iref vdd iref iref iref pfet$5
Xnfet$6_3 vss vss m1_3615_n1223# m1_3615_n1223# m1_3615_n1223# vss nfet$6
Xpfet$5_8 vdd iref vdd iref vdd iref vdd iref iref iref pfet$5
Xpfet$5_9 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$5
.ends

.subckt pfet$8 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
.ends

.subckt nfet$9 a_254_0# a_350_460# a_414_0# a_n84_0# a_94_0# a_510_460# a_190_460#
+ a_574_0# a_30_460# VSUBS
X0 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_460# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_460# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt nfet$7 a_254_0# a_n84_0# a_94_0# a_190_460# a_30_460# VSUBS
X0 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$9 a_254_0# a_348_560# w_n180_n88# a_414_0# a_n92_0# a_94_0# a_574_0#
+ a_508_560# a_188_560# a_28_560#
X0 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt pfet$7 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_348_n136# a_414_0# a_n92_0#
+ a_94_0# a_574_0# a_508_n136#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_n136# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_n136# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$8 a_1054_0# a_734_0# a_254_0# a_350_460# a_830_460# a_894_0# a_990_460#
+ a_1214_0# a_414_0# a_n84_0# a_94_0# a_510_460# a_190_460# a_574_0# a_670_460# a_1150_460#
+ a_30_460# VSUBS
X0 a_734_0# a_670_460# a_574_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_574_0# a_510_460# a_414_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X3 a_1054_0# a_990_460# a_894_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X4 a_894_0# a_830_460# a_734_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X5 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X6 a_414_0# a_350_460# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X7 a_1214_0# a_1150_460# a_1054_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt nfet$10 a_n84_0# a_94_0# a_30_460# VSUBS
X0 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt Ncomparator iref vss vdd inn inp out
Xpfet$8_0 vdd vdd vdd vdd vdd vdd pfet$8
Xpfet$8_1 vdd vdd vdd vdd vdd vdd pfet$8
Xpfet$8_3 vdd vdd vdd vdd vdd vdd pfet$8
Xpfet$8_2 vdd vdd vdd vdd vdd vdd pfet$8
Xnfet$9_0 vss iref m1_506_n191# vss m1_506_n191# iref iref vss iref vss nfet$9
Xnfet$9_1 vss iref iref vss iref iref iref vss iref vss nfet$9
Xnfet$9_2 m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191#
+ m1_506_n191# m1_506_n191# m1_506_n191# vss nfet$9
Xnfet$9_3 m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191#
+ m1_506_n191# m1_506_n191# m1_506_n191# vss nfet$9
Xnfet$7_0 m1_506_n191# m1_506_n191# m1_570_1653# inp inp vss nfet$7
Xnfet$9_5 vss iref m1_506_n191# vss m1_506_n191# iref iref vss iref vss nfet$9
Xnfet$9_4 vss iref iref vss iref iref iref vss iref vss nfet$9
Xnfet$7_1 m1_506_n191# m1_506_n191# m1_1242_549# inn inn vss nfet$7
Xnfet$7_3 m1_506_n191# m1_506_n191# m1_1242_549# inn inn vss nfet$7
Xnfet$7_2 m1_506_n191# m1_506_n191# m1_570_1653# inp inp vss nfet$7
Xpfet$9_0 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$9
Xpfet$9_1 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$9
Xpfet$9_2 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$9
Xpfet$7_0 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_570_1653# vdd m1_570_1653#
+ vdd m1_1242_549# pfet$7
Xpfet$9_3 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$9
Xpfet$7_1 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_1242_549# vdd m1_1242_549#
+ vdd m1_1242_549# pfet$7
Xpfet$7_2 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_570_1653# vdd m1_570_1653#
+ vdd m1_1242_549# pfet$7
Xpfet$7_3 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_1242_549# vdd m1_1242_549#
+ vdd m1_1242_549# pfet$7
Xnfet$8_0 out out vss iref iref vss iref vss out vss out iref iref vss iref iref iref
+ vss nfet$8
Xnfet$10_0 vss vss vss vss nfet$10
Xnfet$10_1 vss vss vss vss nfet$10
.ends

.subckt nfet$11 a_n84_0# a_94_0# a_30_160# VSUBS
X0 a_94_0# a_30_160# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.28u
.ends

.subckt pfet$10 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt SRLATCH vdd vss q qb s r
Xnfet$11_0 vss qb r vss nfet$11
Xnfet$11_1 vss qb q vss nfet$11
Xpfet$10_0 r vdd m1_818_875# qb pfet$10
Xnfet$11_2 q vss s vss nfet$11
Xpfet$10_1 q vdd vdd m1_818_875# pfet$10
Xnfet$11_3 q vss qb vss nfet$11
Xpfet$10_2 s vdd m1_50_875# vdd pfet$10
Xpfet$10_3 qb vdd q m1_50_875# pfet$10
.ends

.subckt ppolyf_u_resistor$2 a_n376_0# a_4200_0# a_n132_0#
X0 a_n132_0# a_4200_0# a_n376_0# ppolyf_u r_width=1u r_length=21u
.ends

.subckt pfet$19 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt pfet$2 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=2.6p pd=9.3u as=2.6p ps=9.3u w=4u l=0.28u
.ends

.subckt nfet$3 a_30_n132# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$3 a_28_460# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_460# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt nfet$2 a_n84_0# a_94_0# a_30_460# VSUBS
X0 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt SCHMITT VDD VSS IN OUT
Xpfet$2_0 IN VDD m1_596_1544# OUT pfet$2
Xpfet$2_1 IN VDD VDD m1_596_1544# pfet$2
Xnfet$3_0 OUT m1_592_402# VDD VSS nfet$3
Xpfet$3_0 OUT VDD m1_596_1544# VSS pfet$3
Xnfet$2_0 m1_592_402# OUT IN VSS nfet$2
Xnfet$2_1 VSS m1_592_402# IN VSS nfet$2
.ends

.subckt VCOfinal_noCP vss vdd irefn qb qnot irefp fout foutb osci
Xnfet$19$1_2 SCHMITT_1/OUT vss fout vss nfet$19$1
Xnfet$19$1_1 SCHMITT_0/OUT vss foutb vss nfet$19$1
XPcomparator_0 vss vdd irefp osci Pcomparator_0/inp SRLATCH_0/r Pcomparator
XNcomparator_0 irefn vss vdd Ncomparator_0/inn osci SRLATCH_0/s Ncomparator
XSRLATCH_0 vdd vss SRLATCH_0/q qb SRLATCH_0/s SRLATCH_0/r SRLATCH
Xppolyf_u_resistor$2_0 vss vss Pcomparator_0/inp ppolyf_u_resistor$2
Xppolyf_u_resistor$2_1 vss m1_13996_n13334# Ncomparator_0/inn ppolyf_u_resistor$2
Xppolyf_u_resistor$2_2 vss m1_13996_n13334# Pcomparator_0/inp ppolyf_u_resistor$2
Xppolyf_u_resistor$2_3 vss vdd Ncomparator_0/inn ppolyf_u_resistor$2
Xpfet$19_0 SRLATCH_0/q vdd vdd qnot pfet$19
Xpfet$19_1 SCHMITT_0/OUT vdd vdd foutb pfet$19
Xpfet$19_2 SCHMITT_1/OUT vdd vdd fout pfet$19
XSCHMITT_0 vdd vss qb SCHMITT_0/OUT SCHMITT
XSCHMITT_1 vdd vss SRLATCH_0/q SCHMITT_1/OUT SCHMITT
Xnfet$19$1_0 SRLATCH_0/q vss qnot vss nfet$19$1
.ends

