* Extracted by KLayout with GF180MCU LVS runset on : 01/09/2025 05:18

.SUBCKT DFF_2phase_1 VSS|VSSd D|Q Q E|PHI_1 D E|PHI_2 VDD|VDDd vss
M$1 VDD|VDDd E|PHI_1 \$2 VDD|VDDd pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$2 \$3 \$2 VDD|VDDd VDD|VDDd pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$3 VDD|VDDd E|PHI_2 \$5 VDD|VDDd pfet_05v0 L=0.5U W=1.38U AS=0.6072P AD=0.476P
+ PS=3.64U PD=2.18U
M$4 \$6 \$5 VDD|VDDd VDD|VDDd pfet_05v0 L=0.5U W=1U AS=0.476P AD=0.44P PS=2.18U
+ PD=2.88U
M$5 \$31 D VDD|VDDd VDD|VDDd pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P PS=2.88U
+ PD=1.24U
M$6 \$10 \$2 \$31 VDD|VDDd pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$7 \$10 \$3 \$32 VDD|VDDd pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$8 VDD|VDDd \$11 \$32 VDD|VDDd pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$9 \$11 \$10 VDD|VDDd VDD|VDDd pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$10 \$37 D|Q VDD|VDDd VDD|VDDd pfet_05v0 L=0.5U W=1U AS=0.44P AD=0.12P
+ PS=2.88U PD=1.24U
M$11 \$13 \$5 \$37 VDD|VDDd pfet_05v0 L=0.5U W=1U AS=0.12P AD=0.26P PS=1.24U
+ PD=1.52U
M$12 \$13 \$6 \$39 VDD|VDDd pfet_05v0 L=0.5U W=1U AS=0.426P AD=0.26P PS=2.08U
+ PD=1.52U
M$13 VDD|VDDd \$14 \$39 VDD|VDDd pfet_05v0 L=0.5U W=1.38U AS=0.426P AD=0.3588P
+ PS=2.08U PD=1.9U
M$14 \$14 \$13 VDD|VDDd VDD|VDDd pfet_05v0 L=0.5U W=1.38U AS=0.3588P AD=0.6072P
+ PS=1.9U PD=3.64U
M$15 VDD|VDDd \$10 D|Q VDD|VDDd pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$16 VDD|VDDd \$13 Q VDD|VDDd pfet_05v0 L=0.5U W=1.83U AS=0.8052P AD=0.8052P
+ PS=4.54U PD=4.54U
M$17 \$18 D VSS|VSSd vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P PS=2.28U
+ PD=0.94U
M$18 \$10 \$3 \$18 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$19 \$19 \$2 \$10 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$20 VSS|VSSd \$11 \$19 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$21 \$11 \$10 VSS|VSSd vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$22 \$25 D|Q VSS|VSSd vss nfet_05v0 L=0.6U W=0.7U AS=0.308P AD=0.084P PS=2.28U
+ PD=0.94U
M$23 \$13 \$6 \$25 vss nfet_05v0 L=0.6U W=0.7U AS=0.084P AD=0.182P PS=0.94U
+ PD=1.22U
M$24 \$21 \$5 \$13 vss nfet_05v0 L=0.6U W=0.7U AS=0.182P AD=0.263P PS=1.22U
+ PD=1.49U
M$25 VSS|VSSd \$14 \$21 vss nfet_05v0 L=0.6U W=0.79U AS=0.263P AD=0.2054P
+ PS=1.49U PD=1.31U
M$26 \$14 \$13 VSS|VSSd vss nfet_05v0 L=0.6U W=0.79U AS=0.2054P AD=0.3476P
+ PS=1.31U PD=2.46U
M$27 VSS|VSSd E|PHI_1 \$2 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$28 \$3 \$2 VSS|VSSd vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$29 VSS|VSSd E|PHI_2 \$5 vss nfet_05v0 L=0.6U W=0.79U AS=0.3476P AD=0.263P
+ PS=2.46U PD=1.49U
M$30 \$6 \$5 VSS|VSSd vss nfet_05v0 L=0.6U W=0.7U AS=0.263P AD=0.308P PS=1.49U
+ PD=2.28U
M$31 VSS|VSSd \$10 D|Q vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
M$32 VSS|VSSd \$13 Q vss nfet_05v0 L=0.6U W=1.32U AS=0.5808P AD=0.5808P
+ PS=3.52U PD=3.52U
.ENDS DFF_2phase_1
