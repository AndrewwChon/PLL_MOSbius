* Extracted by KLayout with GF180MCU LVS runset on : 08/08/2025 05:32

.SUBCKT asc_9_bit_counter A|OUT B|OUT C|OUT D|OUT VSS|vss VDD|vdd E|OUT G|OUT
+ I|OUT F|OUT H|OUT B|Q|clk|in|out B|Q|out A|d1 A|d2 A|d3 A|d4 A|d5 A|d6 A|d7
+ A|d8 A|d9 in|rst clkn|clkp|out ins clkn|clkp|in|out in|ind|ins A|B|out
+ B|ind|ins ins|out OUT|done a|clk|in A|ind|out D|Qb|in vss
M$1 \$12 \$5 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$2 \$13 \$6 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$3 VDD|vdd B|OUT \$5 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$4 \$5 A|OUT VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$5 VDD|vdd \$27 \$6 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$6 \$6 \$12 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$7 \$52 \$24 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$8 \$55 \$14 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$9 \$56 \$16 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$10 \$59 \$17 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$11 \$60 \$25 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$12 \$63 \$19 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$13 \$64 \$21 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$14 \$67 \$22 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$15 \$68 \$26 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$16 \$93 B|Q|clk|in|out A|OUT VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P
+ PS=13.3U PD=13.3U
M$17 \$96 B|Q|clk|in|out B|OUT VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P
+ PS=13.3U PD=13.3U
M$18 \$97 B|Q|clk|in|out C|OUT VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P
+ PS=13.3U PD=13.3U
M$19 \$100 B|Q|clk|in|out D|OUT VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P
+ PS=13.3U PD=13.3U
M$20 \$101 B|Q|clk|in|out E|OUT VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P
+ PS=13.3U PD=13.3U
M$21 \$102 B|Q|clk|in|out F|OUT VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P
+ PS=13.3U PD=13.3U
M$22 \$103 B|Q|clk|in|out G|OUT VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P
+ PS=13.3U PD=13.3U
M$23 \$104 B|Q|clk|in|out H|OUT VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P
+ PS=13.3U PD=13.3U
M$24 \$105 B|Q|out I|OUT VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$25 VDD|vdd A|d1 \$93 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$26 VDD|vdd A|d2 \$96 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$27 VDD|vdd A|d3 \$97 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$28 VDD|vdd A|d4 \$100 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$29 VDD|vdd A|d5 \$101 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$30 VDD|vdd A|d6 \$102 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$31 VDD|vdd A|d7 \$103 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$32 VDD|vdd A|d8 \$104 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$33 VDD|vdd A|d9 \$105 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$34 A|OUT \$180 \$52 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$35 B|OUT \$181 \$55 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$36 C|OUT \$182 \$56 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$37 D|OUT \$183 \$59 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$38 E|OUT \$184 \$60 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$39 F|OUT \$185 \$63 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$40 G|OUT \$186 \$64 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$41 H|OUT \$187 \$67 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$42 I|OUT \$188 \$68 VDD|vdd pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U
+ PD=13.3U
M$43 VDD|vdd C|OUT \$155 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$44 \$155 D|OUT VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$45 \$27 \$155 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$46 VDD|vdd \$13 \$157 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$47 \$157 \$247 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$48 \$149 \$157 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$49 \$180 B|Q|clk|in|out VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$50 \$24 A|d1 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$51 VDD|vdd A|d2 \$14 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$52 VDD|vdd B|Q|clk|in|out \$181 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$53 \$182 B|Q|clk|in|out VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$54 \$16 A|d3 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$55 VDD|vdd A|d4 \$17 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$56 VDD|vdd B|Q|clk|in|out \$183 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$57 \$184 B|Q|clk|in|out VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$58 \$25 A|d5 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$59 VDD|vdd A|d6 \$19 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$60 VDD|vdd B|Q|clk|in|out \$185 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$61 \$186 B|Q|clk|in|out VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$62 \$21 A|d7 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$63 VDD|vdd A|d8 \$22 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$64 VDD|vdd B|Q|clk|in|out \$187 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$65 \$188 B|Q|out VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$66 \$26 A|d9 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$67 clkn|clkp|in|out a|clk|in VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$68 clkn|clkp|out clkn|clkp|in|out VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=27U
+ AS=17.55P AD=17.55P PS=65.7U PD=65.7U
M$69 VDD|vdd A|ind|out ins VDD|vdd pfet_03v3 L=0.5U W=27U AS=17.55P AD=17.55P
+ PS=65.7U PD=65.7U
M$70 ins A|B|out VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=27U AS=17.55P AD=17.55P
+ PS=65.7U PD=65.7U
M$71 VDD|vdd in|rst A|B|out VDD|vdd pfet_03v3 L=0.5U W=27U AS=17.55P AD=17.55P
+ PS=65.7U PD=65.7U
M$72 VDD|vdd D|Qb|in ins|out VDD|vdd pfet_03v3 L=0.5U W=27U AS=17.55P AD=17.55P
+ PS=65.7U PD=65.7U
M$73 clkn|clkp|in|out B|Q|clk|in|out VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=24U
+ AS=15.6P AD=15.6P PS=58.4U PD=58.4U
M$83 VDD|vdd F|OUT \$358 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$84 \$358 E|OUT VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$85 \$438 \$358 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$86 VDD|vdd I|OUT \$360 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$87 \$360 \$149 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$88 OUT|done \$360 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$89 ins clkn|clkp|in|out in|ind|ins VDD|vdd pfet_03v3 L=0.5U W=27U AS=17.55P
+ AD=17.55P PS=65.7U PD=65.7U
M$90 ins|out clkn|clkp|out B|ind|ins VDD|vdd pfet_03v3 L=0.5U W=27U AS=17.55P
+ AD=17.55P PS=65.7U PD=65.7U
M$105 VDD|vdd G|OUT \$506 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$106 \$506 H|OUT VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$107 VDD|vdd \$438 \$508 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$108 \$508 \$573 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$109 in|ind|ins clkn|clkp|out \$590 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$110 B|ind|ins clkn|clkp|in|out A|ind|out VDD|vdd pfet_03v3 L=0.5U W=27U
+ AS=17.55P AD=17.55P PS=65.7U PD=65.7U
M$111 in|ind|ins clkn|clkp|out \$591 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$113 \$573 \$506 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$114 \$247 \$508 VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$115 in|ind|ins clkn|clkp|out \$592 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$117 in|ind|ins clkn|clkp|out \$593 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$119 \$590 D|Qb|in VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$120 A|ind|out in|ind|ins VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=27U AS=17.55P
+ AD=17.55P PS=65.7U PD=65.7U
M$121 B|Q|clk|in|out D|Qb|in VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=24U AS=15.6P
+ AD=15.6P PS=58.4U PD=58.4U
M$122 \$591 D|Qb|in VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$125 \$592 D|Qb|in VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$127 \$593 D|Qb|in VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$129 VDD|vdd A|B|out D|Qb|in VDD|vdd pfet_03v3 L=0.5U W=27U AS=17.55P
+ AD=17.55P PS=65.7U PD=65.7U
M$130 D|Qb|in B|ind|ins VDD|vdd VDD|vdd pfet_03v3 L=0.5U W=27U AS=17.55P
+ AD=17.55P PS=65.7U PD=65.7U
M$149 VDD|vdd D|Qb|in B|Q|out VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$151 VDD|vdd D|Qb|in \$749 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$154 VDD|vdd D|Qb|in \$754 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$157 VDD|vdd D|Qb|in \$759 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$160 VDD|vdd D|Qb|in \$764 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$163 VDD|vdd D|Qb|in \$769 VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$169 \$749 clkn|clkp|out in|ind|ins VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$177 \$754 clkn|clkp|out in|ind|ins VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$183 \$759 clkn|clkp|out in|ind|ins VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$187 \$764 clkn|clkp|out in|ind|ins VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$191 \$769 clkn|clkp|out in|ind|ins VDD|vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$214 \$53 \$24 A|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$215 \$54 \$14 B|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$216 \$57 \$16 C|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$217 \$58 \$17 D|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$218 \$61 \$25 E|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$219 \$62 \$19 F|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$220 \$65 \$21 G|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$221 \$66 \$22 H|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$222 \$69 \$26 I|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$223 VSS|vss B|Q|clk|in|out \$53 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$224 VSS|vss B|Q|clk|in|out \$54 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$225 VSS|vss B|Q|clk|in|out \$57 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$226 VSS|vss B|Q|clk|in|out \$58 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$227 VSS|vss B|Q|clk|in|out \$61 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$228 VSS|vss B|Q|clk|in|out \$62 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$229 VSS|vss B|Q|clk|in|out \$65 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$230 VSS|vss B|Q|clk|in|out \$66 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$231 VSS|vss B|Q|out \$69 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$232 \$12 \$5 VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$233 \$13 \$6 VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$234 \$109 B|OUT VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$235 \$5 A|OUT \$109 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$236 \$110 \$27 VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$237 \$6 \$12 \$110 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$238 \$132 A|d1 A|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$239 \$133 A|d2 B|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$240 \$136 A|d3 C|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$241 \$137 A|d4 D|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$242 \$140 A|d5 E|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$243 \$141 A|d6 F|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$244 \$144 A|d7 G|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$245 \$145 A|d8 H|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$246 \$148 A|d9 I|OUT vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$247 \$27 \$155 VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$248 \$149 \$157 VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$249 VSS|vss \$180 \$132 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$250 VSS|vss \$181 \$133 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$251 VSS|vss \$182 \$136 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$252 VSS|vss \$183 \$137 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$253 VSS|vss \$184 \$140 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$254 VSS|vss \$185 \$141 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$255 VSS|vss \$186 \$144 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$256 VSS|vss \$187 \$145 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$257 VSS|vss \$188 \$148 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$258 \$180 B|Q|clk|in|out VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$259 \$24 A|d1 VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$260 VSS|vss A|d2 \$14 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$261 VSS|vss B|Q|clk|in|out \$181 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$262 \$182 B|Q|clk|in|out VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$263 \$16 A|d3 VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$264 VSS|vss A|d4 \$17 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$265 VSS|vss B|Q|clk|in|out \$183 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$266 \$184 B|Q|clk|in|out VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$267 \$25 A|d5 VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$268 VSS|vss A|d6 \$19 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$269 VSS|vss B|Q|clk|in|out \$185 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$270 \$186 B|Q|clk|in|out VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$271 \$21 A|d7 VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$272 VSS|vss A|d8 \$22 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$273 VSS|vss B|Q|clk|in|out \$187 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$274 \$188 B|Q|out VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$275 \$26 A|d9 VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$276 \$191 C|OUT VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$277 \$155 D|OUT \$191 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$278 \$192 \$13 VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$279 \$157 \$247 \$192 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$280 clkn|clkp|in|out a|clk|in VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P
+ AD=0.61P PS=3.22U PD=3.22U
M$281 clkn|clkp|out clkn|clkp|in|out VSS|vss vss nfet_03v3 L=0.5U W=9U AS=5.49P
+ AD=5.49P PS=28.98U PD=28.98U
M$282 ins clkn|clkp|out in|ind|ins vss nfet_03v3 L=0.5U W=9U AS=5.49P AD=5.49P
+ PS=28.98U PD=28.98U
M$283 VSS|vss in|rst A|B|out vss nfet_03v3 L=0.5U W=9U AS=5.49P AD=5.49P
+ PS=28.98U PD=28.98U
M$284 ins|out clkn|clkp|in|out B|ind|ins vss nfet_03v3 L=0.5U W=9U AS=5.49P
+ AD=5.49P PS=28.98U PD=28.98U
M$285 VSS|vss D|Qb|in ins|out vss nfet_03v3 L=0.5U W=9U AS=5.49P AD=5.49P
+ PS=28.98U PD=28.98U
M$286 clkn|clkp|in|out B|Q|clk|in|out VSS|vss vss nfet_03v3 L=0.5U W=8U
+ AS=4.88P AD=4.88P PS=25.76U PD=25.76U
M$296 \$450 F|OUT VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$297 \$358 E|OUT \$450 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$298 \$438 \$358 VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$299 \$451 I|OUT VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$300 \$360 \$149 \$451 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$301 OUT|done \$360 VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$302 \$501 A|ind|out ins vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$303 VSS|vss A|B|out \$501 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$304 \$502 A|ind|out ins vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$305 VSS|vss A|B|out \$502 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$308 \$503 A|ind|out ins vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$309 VSS|vss A|B|out \$503 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$314 \$504 A|ind|out ins vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$315 VSS|vss A|B|out \$504 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$318 \$505 G|OUT VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$319 \$506 H|OUT \$505 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$320 \$507 \$438 VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$321 \$508 \$573 \$507 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$322 \$590 D|Qb|in VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$323 in|ind|ins clkn|clkp|in|out \$590 vss nfet_03v3 L=0.5U W=1U AS=0.61P
+ AD=0.61P PS=3.22U PD=3.22U
M$324 A|ind|out in|ind|ins VSS|vss vss nfet_03v3 L=0.5U W=9U AS=5.49P AD=5.49P
+ PS=28.98U PD=28.98U
M$325 A|ind|out clkn|clkp|out B|ind|ins vss nfet_03v3 L=0.5U W=9U AS=5.49P
+ AD=5.49P PS=28.98U PD=28.98U
M$327 \$586 B|ind|ins VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$328 D|Qb|in A|B|out \$586 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$329 \$749 clkn|clkp|in|out in|ind|ins vss nfet_03v3 L=0.5U W=1U AS=0.61P
+ AD=0.61P PS=3.22U PD=3.22U
M$330 B|Q|clk|in|out D|Qb|in VSS|vss vss nfet_03v3 L=0.5U W=8U AS=4.88P
+ AD=4.88P PS=25.76U PD=25.76U
M$331 \$591 D|Qb|in VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$332 in|ind|ins clkn|clkp|in|out \$591 vss nfet_03v3 L=0.5U W=1U AS=0.61P
+ AD=0.61P PS=3.22U PD=3.22U
M$336 \$587 B|ind|ins VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$337 D|Qb|in A|B|out \$587 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$338 \$754 clkn|clkp|in|out in|ind|ins vss nfet_03v3 L=0.5U W=1U AS=0.61P
+ AD=0.61P PS=3.22U PD=3.22U
M$340 \$592 D|Qb|in VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$341 in|ind|ins clkn|clkp|in|out \$592 vss nfet_03v3 L=0.5U W=1U AS=0.61P
+ AD=0.61P PS=3.22U PD=3.22U
M$345 \$588 B|ind|ins VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$346 D|Qb|in A|B|out \$588 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$347 \$759 clkn|clkp|in|out in|ind|ins vss nfet_03v3 L=0.5U W=1U AS=0.61P
+ AD=0.61P PS=3.22U PD=3.22U
M$349 \$593 D|Qb|in VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$350 in|ind|ins clkn|clkp|in|out \$593 vss nfet_03v3 L=0.5U W=1U AS=0.61P
+ AD=0.61P PS=3.22U PD=3.22U
M$354 \$589 B|ind|ins VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$355 D|Qb|in A|B|out \$589 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$356 \$764 clkn|clkp|in|out in|ind|ins vss nfet_03v3 L=0.5U W=1U AS=0.61P
+ AD=0.61P PS=3.22U PD=3.22U
M$359 \$769 clkn|clkp|in|out in|ind|ins vss nfet_03v3 L=0.5U W=1U AS=0.61P
+ AD=0.61P PS=3.22U PD=3.22U
M$360 \$573 \$506 VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$361 \$247 \$508 VSS|vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$362 VSS|vss D|Qb|in B|Q|out vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$364 VSS|vss D|Qb|in \$749 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$367 VSS|vss D|Qb|in \$754 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$370 VSS|vss D|Qb|in \$759 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$373 VSS|vss D|Qb|in \$764 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$376 VSS|vss D|Qb|in \$769 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$378 \$821 A|B|out D|Qb|in vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$379 VSS|vss B|ind|ins \$821 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$381 \$896 A|B|out VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$382 ins A|ind|out \$896 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$386 \$823 A|B|out D|Qb|in vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$387 VSS|vss B|ind|ins \$823 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$389 \$898 A|B|out VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$390 ins A|ind|out \$898 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$393 \$825 A|B|out D|Qb|in vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$394 VSS|vss B|ind|ins \$825 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$395 \$900 A|B|out VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$396 ins A|ind|out \$900 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$397 \$827 A|B|out D|Qb|in vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$398 VSS|vss B|ind|ins \$827 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$399 \$902 A|B|out VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$400 ins A|ind|out \$902 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$401 \$829 A|B|out D|Qb|in vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$402 VSS|vss B|ind|ins \$829 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$403 \$904 A|B|out VSS|vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P
+ PS=5.22U PD=5.22U
M$404 ins A|ind|out \$904 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
.ENDS asc_9_bit_counter
