** sch_path: /foss/designs/libs/core_analog/asc_hysteresis_buffer/asc_hysteresis_buffer.sch
.subckt asc_hysteresis_buffer in vss out vdd
*.PININFO in:B out:B vss:B vdd:B
M1 net1 in vdd vdd pfet_03v3 L=0.5u W=3.0u nf=1 m=1
M2 net1 in vss vss nfet_03v3 L=0.5u W=1.0u nf=1 m=1
M3 net2 net1 vdd vdd pfet_03v3 L=0.5u W=12.0u nf=1 m=1
M4 net2 net1 vss vss nfet_03v3 L=0.5u W=4.0u nf=1 m=1
M5 net3 net2 vdd vdd pfet_03v3 L=0.5u W=48.0u nf=4 m=1
M6 net3 net2 vss vss nfet_03v3 L=0.5u W=16.0u nf=4 m=1
M7 out net3 vdd vdd pfet_03v3 L=0.5u W=96.0u nf=8 m=1
M8 out net3 vss vss nfet_03v3 L=0.5u W=32.0u nf=8 m=1
x1 net3 vdd net2 vss inv1u05u
.ends

* expanding   symbol:  libs/core_analog/inv1u05u/inv1u05u.sym # of pins=4
** sym_path: /foss/designs/libs/core_analog/inv1u05u/inv1u05u.sym
** sch_path: /foss/designs/libs/core_analog/inv1u05u/inv1u05u.sch
.subckt inv1u05u in vdd out vss
*.PININFO in:B out:B vss:B vdd:B
M1 out in vdd vdd pfet_03v3 L=0.5u W=3.0u nf=1 m=1
M2 out in vss vss nfet_03v3 L=0.5u W=1.0u nf=1 m=1
.ends

