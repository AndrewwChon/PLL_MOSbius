* Extracted by KLayout with GF180MCU LVS runset on : 07/08/2025 03:22

.SUBCKT asc_SR_ltch
M$1 \$15 S VDD VDD pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U PD=13.3U
M$2 Qb Q \$15 VDD pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U PD=13.3U
M$3 \$16 R VDD VDD pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U PD=13.3U
M$4 Q Qb \$16 VDD pfet_03v3 L=0.5U W=6U AS=3.9P AD=3.9P PS=13.3U PD=13.3U
M$5 Qb S VSS VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$6 VSS Q Qb VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$7 Q R VSS VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$8 VSS Qb Q VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
.ENDS asc_SR_ltch
