** sch_path: /foss/designs/libs/core_analog/asc_mim_cap_lvs_test/asc_mim_cap_lvs_test.sch
.subckt asc_mim_cap_lvs_test vin vss
*.PININFO vin:B vss:B
XM1 net2 vin net1 vss nfet_03v3 L=0.5u W=1u nf=1 m=1
XC2 net1 vss cap_mim_2f0fF c_width=10e-6 c_length=5e-6 m=1
XC4 net2 vss cap_mim_2f0fF c_width=10e-6 c_length=5e-6 m=1
.ends
