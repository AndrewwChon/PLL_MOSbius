* Extracted by KLayout with GF180MCU LVS runset on : 13/08/2025 22:03

.SUBCKT xp_programmable_basic_pump vss out down iref vdd s1 s2 s3 s4 up
M$1 vdd s1 \$30 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$2 vdd s2 \$36 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$3 vdd s3 \$38 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$4 vdd s4 \$40 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$5 vdd up \$127 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$6 \$94 \$30 \$34 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$7 iref \$30 \$54 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$8 \$94 s1 vdd vdd pfet_03v3 L=0.5U W=1U AS=0.65P AD=0.65P PS=3.3U PD=3.3U
M$9 \$95 \$36 \$34 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$10 iref \$36 \$23 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$11 \$95 s2 vdd vdd pfet_03v3 L=0.5U W=1U AS=0.65P AD=0.65P PS=3.3U PD=3.3U
M$12 \$96 \$38 \$34 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$13 iref \$38 \$4 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$14 \$96 s3 vdd vdd pfet_03v3 L=0.5U W=1U AS=0.65P AD=0.65P PS=3.3U PD=3.3U
M$15 \$126 \$40 \$34 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$16 iref \$40 \$8 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$17 \$126 s4 vdd vdd pfet_03v3 L=0.5U W=1U AS=0.65P AD=0.65P PS=3.3U PD=3.3U
M$18 vdd vdd vdd vdd pfet_03v3 L=0.5U W=168U AS=94.71P AD=94.71P PS=300.06U
+ PD=300.06U
M$19 out \$126 \$128 vdd pfet_03v3 L=0.5U W=336U AS=109.2P AD=109.2P PS=423.2U
+ PD=423.2U
M$31 out \$96 \$125 vdd pfet_03v3 L=0.5U W=168U AS=54.6P AD=54.6P PS=211.6U
+ PD=211.6U
M$57 \$128 \$127 vdd vdd pfet_03v3 L=0.5U W=336U AS=96.32P AD=96.32P PS=363.52U
+ PD=363.52U
M$69 \$125 \$127 vdd vdd pfet_03v3 L=0.5U W=168U AS=48.16P AD=48.16P PS=181.76U
+ PD=181.76U
M$98 out \$95 \$140 vdd pfet_03v3 L=0.5U W=84U AS=27.3P AD=27.3P PS=105.8U
+ PD=105.8U
M$104 out \$94 \$142 vdd pfet_03v3 L=0.5U W=42U AS=13.65P AD=13.65P PS=52.9U
+ PD=52.9U
M$110 \$34 \$34 \$141 vdd pfet_03v3 L=0.5U W=42U AS=13.65P AD=13.65P PS=52.9U
+ PD=52.9U
M$168 \$140 \$127 vdd vdd pfet_03v3 L=0.5U W=84U AS=24.08P AD=24.08P PS=90.88U
+ PD=90.88U
M$174 \$142 \$127 vdd vdd pfet_03v3 L=0.5U W=42U AS=12.04P AD=12.04P PS=45.44U
+ PD=45.44U
M$180 \$141 vss vdd vdd pfet_03v3 L=0.5U W=42U AS=12.04P AD=12.04P PS=45.44U
+ PD=45.44U
M$234 vss vss vss vss nfet_03v3 L=0.5U W=168U AS=68.67P AD=68.67P PS=250.62U
+ PD=250.62U
M$236 out \$8 \$17 vss nfet_03v3 L=0.5U W=112U AS=48.72P AD=48.72P PS=181.92U
+ PD=181.92U
M$240 out \$4 \$5 vss nfet_03v3 L=0.5U W=56U AS=24.36P AD=24.36P PS=90.96U
+ PD=90.96U
M$252 \$17 down vss vss nfet_03v3 L=0.5U W=112U AS=36.96P AD=36.96P PS=122.56U
+ PD=122.56U
M$256 \$5 down vss vss nfet_03v3 L=0.5U W=56U AS=18.48P AD=18.48P PS=61.28U
+ PD=61.28U
M$268 \$20 down vss vss nfet_03v3 L=0.5U W=28U AS=9.24P AD=9.24P PS=30.64U
+ PD=30.64U
M$270 \$31 vdd vss vss nfet_03v3 L=0.5U W=14U AS=4.62P AD=4.62P PS=15.32U
+ PD=15.32U
M$272 \$32 down vss vss nfet_03v3 L=0.5U W=14U AS=4.62P AD=4.62P PS=15.32U
+ PD=15.32U
M$274 \$33 vdd vss vss nfet_03v3 L=0.5U W=14U AS=4.62P AD=4.62P PS=15.32U
+ PD=15.32U
M$282 out \$23 \$20 vss nfet_03v3 L=0.5U W=28U AS=12.18P AD=12.18P PS=45.48U
+ PD=45.48U
M$284 iref iref \$31 vss nfet_03v3 L=0.5U W=14U AS=6.09P AD=6.09P PS=22.74U
+ PD=22.74U
M$286 out \$54 \$32 vss nfet_03v3 L=0.5U W=14U AS=6.09P AD=6.09P PS=22.74U
+ PD=22.74U
M$288 \$34 iref \$33 vss nfet_03v3 L=0.5U W=14U AS=6.09P AD=6.09P PS=22.74U
+ PD=22.74U
M$310 vss \$30 \$54 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$311 vss s1 \$30 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$312 iref s1 \$54 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$313 vss \$36 \$23 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$314 iref s2 \$23 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$315 vss s2 \$36 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$316 vss \$38 \$4 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$317 vss s3 \$38 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$318 iref s3 \$4 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$319 vss \$40 \$8 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$320 iref s4 \$8 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$321 vss s4 \$40 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$322 vss up \$127 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$339 \$94 s1 \$34 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$340 \$95 s2 \$34 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$341 \$96 s3 \$34 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$342 \$126 s4 \$34 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
.ENDS xp_programmable_basic_pump
