* Extracted by KLayout with GF180MCU LVS runset on : 12/08/2025 07:07

.SUBCKT PLAY D|VSS G VSS
M$1 \$3 G D|VSS VSS nfet_03v3 L=0.5U W=14U AS=6.09P AD=6.09P PS=22.74U PD=22.74U
M$3 D|VSS G D|VSS VSS nfet_03v3 L=0.5U W=14U AS=6.09P AD=6.09P PS=22.74U
+ PD=22.74U
.ENDS PLAY
