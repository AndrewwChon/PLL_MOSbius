* NGSPICE file created from scan_chain.ext - technology: gf180mcuD

.subckt nfet$2 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt pfet$2 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$3 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$1 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt nfet a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt pfet$3 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$1 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt qw_NOLclk CLK VDDd VSSd PHI_2 PHI_1
Xnfet$2_2 m1_11601_2380# VSSd PHI_2 VSSd nfet$2
Xpfet_0 VDDd VDDd m1_13930_233# PHI_1 pfet
Xpfet_1 VDDd VDDd m1_13930_1818# PHI_2 pfet
Xnfet$2_3 CLK VSSd m1_11161_409# VSSd nfet$2
Xpfet$2_0 VDDd VDDd PHI_1 m1_11601_71# pfet$2
Xpfet$2_1 VDDd VDDd m1_11379_n171# m1_11161_409# pfet$2
Xpfet$2_2 VDDd VDDd PHI_2 m1_11601_2380# pfet$2
Xpfet$2_3 VDDd VDDd m1_11161_409# CLK pfet$2
Xnfet$3_0 m1_12351_431# m1_12351_431# m1_11601_71# m1_11601_71# m1_11837_749# VSSd
+ nfet$3
Xnfet$3_1 m1_11379_n171# m1_11379_n171# VSSd VSSd m1_11837_749# VSSd nfet$3
Xnfet$3_2 m1_12351_2064# m1_12351_2064# m1_11601_2380# m1_11601_2380# m1_11837_1708#
+ VSSd nfet$3
Xnfet$3_3 m1_11161_409# m1_11161_409# VSSd VSSd m1_11837_1708# VSSd nfet$3
Xnfet$1_0 m1_12351_2064# m1_15103_233# VSSd VSSd nfet$1
Xnfet$1_1 m1_15103_233# m1_13930_233# VSSd VSSd nfet$1
Xnfet$1_2 m1_12351_431# m1_15103_1818# VSSd VSSd nfet$1
Xnfet$1_3 m1_15103_1818# m1_13930_1818# VSSd VSSd nfet$1
Xnfet_0 PHI_1 VSSd m1_13930_233# VSSd nfet
Xnfet_1 PHI_2 VSSd m1_13930_1818# VSSd nfet
Xpfet$3_0 VDDd m1_11601_71# VDDd m1_11379_n171# pfet$3
Xpfet$3_1 VDDd VDDd m1_11601_71# m1_12351_431# pfet$3
Xpfet$3_2 VDDd m1_11601_2380# VDDd m1_11161_409# pfet$3
Xpfet$3_3 VDDd VDDd m1_11601_2380# m1_12351_2064# pfet$3
Xpfet$1_0 m1_12351_2064# VDDd VDDd m1_15103_233# pfet$1
Xpfet$1_1 m1_15103_233# VDDd VDDd m1_13930_233# pfet$1
Xpfet$1_2 m1_12351_431# VDDd VDDd m1_15103_1818# pfet$1
Xpfet$1_3 m1_15103_1818# VDDd VDDd m1_13930_1818# pfet$1
Xnfet$2_0 m1_11601_71# VSSd PHI_1 VSSd nfet$2
Xnfet$2_1 m1_11161_409# VSSd m1_11379_n171# VSSd nfet$2
.ends

.subckt pfet$8 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$6 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$9 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$7 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$10 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$9 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$7 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$8 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$6 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$10 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_hysteresis_buffer vss in vdd out
Xpfet$8_0 vdd vdd m1_348_648# in pfet$8
Xpfet$6_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd m1_884_42#
+ m1_884_42# pfet$6
Xnfet$9_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$9
Xnfet$7_0 m1_348_648# vss m1_884_42# vss nfet$7
Xpfet$10_0 vdd vdd m1_884_42# m1_1156_42# pfet$10
Xpfet$9_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$9
Xpfet$7_0 vdd vdd m1_884_42# m1_348_648# pfet$7
Xnfet$8_0 in vss m1_348_648# vss nfet$8
Xnfet$6_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$6
Xnfet$10_0 m1_1156_42# vss m1_884_42# vss nfet$10
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__latq_1$2 D E Q VDD VSS VNW VPW
X0 VSS a_1020_652# Q VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X1 a_504_110# a_36_92# VDD VNW pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X2 VDD a_1020_652# Q VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X3 a_1264_107# a_36_92# a_1020_652# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X4 VSS E a_36_92# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X5 VSS a_1364_532# a_1264_107# VPW nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X6 VDD E a_36_92# VNW pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X7 VDD a_1364_532# a_1224_652# VNW pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X8 a_872_652# D VDD VNW pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X9 a_1364_532# a_1020_652# VDD VNW pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X10 a_1020_652# a_504_110# a_872_107# VPW nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X11 a_872_107# D VSS VPW nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X12 a_1020_652# a_36_92# a_872_652# VNW pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X13 a_504_110# a_36_92# VSS VPW nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X14 a_1364_532# a_1020_652# VSS VPW nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X15 a_1224_652# a_504_110# a_1020_652# VNW pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt DFF_2phase_1$1 D PHI_2 PHI_1 Q VDDd VSSd
Xgf180mcu_fd_sc_mcu9t5v0__latq_1$2_0 gf180mcu_fd_sc_mcu9t5v0__latq_1$2_1/Q PHI_2 Q
+ VDDd VSSd VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1$2
Xgf180mcu_fd_sc_mcu9t5v0__latq_1$2_1 D PHI_1 gf180mcu_fd_sc_mcu9t5v0__latq_1$2_1/Q
+ VDDd VSSd VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1$2
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1$1 I VDD VSS ZN VNW VPW
X0 ZN I VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__and2_1$1 A1 A2 VDD VSS Z VNW VPW
X0 VDD A2 a_36_201# VNW pfet_05v0 ad=0.5054p pd=2.57u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1 a_244_201# A1 a_36_201# VPW nfet_05v0 ad=0.1056p pd=0.98u as=0.2904p ps=2.2u w=0.66u l=0.6u
X2 Z a_36_201# VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.3894p ps=2.06u w=1.32u l=0.6u
X3 Z a_36_201# VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.5054p ps=2.57u w=1.83u l=0.5u
X4 VSS A2 a_244_201# VPW nfet_05v0 ad=0.3894p pd=2.06u as=0.1056p ps=0.98u w=0.66u l=0.6u
X5 a_36_201# A1 VDD VNW pfet_05v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__or2_1$1 A1 A2 VDD VSS Z VNW VPW
X0 a_255_756# A1 a_67_756# VNW pfet_05v0 ad=0.2379p pd=1.435u as=0.4026p ps=2.71u w=0.915u l=0.5u
X1 VSS A2 a_67_756# VPW nfet_05v0 ad=0.3828p pd=2.08u as=0.1716p ps=1.18u w=0.66u l=0.6u
X2 VDD A2 a_255_756# VNW pfet_05v0 ad=0.57645p pd=2.69u as=0.2379p ps=1.435u w=0.915u l=0.5u
X3 Z a_67_756# VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.3828p ps=2.08u w=1.32u l=0.6u
X4 Z a_67_756# VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.57645p ps=2.69u w=1.83u l=0.5u
X5 a_67_756# A1 VSS VPW nfet_05v0 ad=0.1716p pd=1.18u as=0.2904p ps=2.2u w=0.66u l=0.6u
.ends

.subckt Register_unitcell out q default phi2 phi1 en d VSSd VDDd
XDFF_2phase_1$1_0 d phi2 phi1 q VDDd VSSd DFF_2phase_1$1
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$1_0 en VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1$1
Xgf180mcu_fd_sc_mcu9t5v0__and2_1$1_0 gf180mcu_fd_sc_mcu9t5v0__inv_1$1_0/ZN default
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1$1_0/A1 VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1$1
Xgf180mcu_fd_sc_mcu9t5v0__and2_1$1_1 q en VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1$1_0/A2
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1$1
Xgf180mcu_fd_sc_mcu9t5v0__or2_1$1_0 gf180mcu_fd_sc_mcu9t5v0__or2_1$1_0/A1 gf180mcu_fd_sc_mcu9t5v0__or2_1$1_0/A2
+ VDDd VSSd out VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1$1
.ends

.subckt SRegister_10$1 out[1] out[2] out[3] out[9] d q default10 default9 default8
+ default7 default6 default5 default4 default3 default2 default1 out[6] out[4] out[10]
+ out[7] out[5] out[8] phi2 en VDDd phi1 VSSd
XRegister_unitcell_0 out[2] Register_unitcell_7/d default2 phi2 phi1 en Register_unitcell_6/q
+ VSSd VDDd Register_unitcell
XRegister_unitcell_1 out[6] Register_unitcell_2/d default6 phi2 phi1 en Register_unitcell_9/q
+ VSSd VDDd Register_unitcell
XRegister_unitcell_2 out[7] Register_unitcell_3/d default7 phi2 phi1 en Register_unitcell_2/d
+ VSSd VDDd Register_unitcell
XRegister_unitcell_3 out[8] Register_unitcell_4/d default8 phi2 phi1 en Register_unitcell_3/d
+ VSSd VDDd Register_unitcell
XRegister_unitcell_5 out[10] q default10 phi2 phi1 en Register_unitcell_5/d VSSd VDDd
+ Register_unitcell
XRegister_unitcell_4 out[9] Register_unitcell_5/d default9 phi2 phi1 en Register_unitcell_4/d
+ VSSd VDDd Register_unitcell
XRegister_unitcell_6 out[1] Register_unitcell_6/q default1 phi2 phi1 en d VSSd VDDd
+ Register_unitcell
XRegister_unitcell_7 out[3] Register_unitcell_8/d default3 phi2 phi1 en Register_unitcell_7/d
+ VSSd VDDd Register_unitcell
XRegister_unitcell_8 out[4] Register_unitcell_9/d default4 phi2 phi1 en Register_unitcell_8/d
+ VSSd VDDd Register_unitcell
XRegister_unitcell_9 out[5] Register_unitcell_9/q default5 phi2 phi1 en Register_unitcell_9/d
+ VSSd VDDd Register_unitcell
.ends

.subckt pfet$4 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=2.6p pd=9.3u as=2.6p ps=9.3u w=4u l=0.28u
.ends

.subckt nfet$5 a_30_n132# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$5 a_28_460# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_460# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt nfet$4 a_n84_0# a_94_0# a_30_460# VSUBS
X0 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt SCHMITT VDD VSS IN OUT
Xpfet$4_0 IN VDD m1_596_1544# OUT pfet$4
Xpfet$4_1 IN VDD VDD m1_596_1544# pfet$4
Xnfet$5_0 OUT m1_592_402# VDD VSS nfet$5
Xpfet$5_0 OUT VDD m1_596_1544# VSS pfet$5
Xnfet$4_0 m1_592_402# OUT IN VSS nfet$4
Xnfet$4_1 VSS m1_592_402# IN VSS nfet$4
.ends

.subckt scan_chain VDDd VSSd ENd DATAd CLKd out[1] out[2] out[3] out[4] out[5] out[6]
+ out[7] out[8] out[9] out[10] out[20] out[19] out[18] out[17] out[16] out[15] out[14]
+ out[13] out[12] out[11] out[21] out[22] out[23] out[24] out[25] out[26] out[27]
+ out[28] out[29] out[30] out[40] out[39] out[38] out[37] out[36] out[35] out[34]
+ out[33] out[32] out[31] out[41] out[42] out[43] out[44] out[45] out[46] out[47]
+ out[48] out[49] out[50]
Xqw_NOLclk_0 SCHMITT_0/OUT VDDd VSSd qw_NOLclk_0/PHI_2 qw_NOLclk_0/PHI_1 qw_NOLclk
Xasc_hysteresis_buffer_0 VSSd CLKd VDDd SCHMITT_0/IN asc_hysteresis_buffer
XSRegister_10$1_0 out[31] out[32] out[33] out[39] SRegister_10$1_3/q SRegister_10$1_2/d
+ VSSd VSSd VDDd VSSd VSSd VDDd VDDd VSSd VSSd VSSd out[36] out[34] out[40] out[37]
+ out[35] out[38] qw_NOLclk_0/PHI_2 SRegister_10$1_4/en VDDd qw_NOLclk_0/PHI_1 VSSd
+ SRegister_10$1
Xasc_hysteresis_buffer_1 VSSd ENd VDDd SRegister_10$1_4/en asc_hysteresis_buffer
XSRegister_10$1_1 out[11] out[12] out[13] out[19] SRegister_10$1_4/q SRegister_10$1_3/d
+ VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd out[16] out[14] out[20] out[17]
+ out[15] out[18] qw_NOLclk_0/PHI_2 SRegister_10$1_4/en VDDd qw_NOLclk_0/PHI_1 VSSd
+ SRegister_10$1
Xasc_hysteresis_buffer_2 VSSd DATAd VDDd SRegister_10$1_4/d asc_hysteresis_buffer
XSRegister_10$1_2 out[41] out[42] out[43] out[49] SRegister_10$1_2/d SRegister_10$1_2/q
+ VSSd VSSd VSSd VSSd VDDd VSSd VSSd VDDd VDDd VSSd out[46] out[44] out[50] out[47]
+ out[45] out[48] qw_NOLclk_0/PHI_2 SRegister_10$1_4/en VDDd qw_NOLclk_0/PHI_1 VSSd
+ SRegister_10$1
XSRegister_10$1_3 out[21] out[22] out[23] out[29] SRegister_10$1_3/d SRegister_10$1_3/q
+ VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd out[26] out[24] out[30] out[27]
+ out[25] out[28] qw_NOLclk_0/PHI_2 SRegister_10$1_4/en VDDd qw_NOLclk_0/PHI_1 VSSd
+ SRegister_10$1
XSRegister_10$1_4 out[1] out[2] out[3] out[9] SRegister_10$1_4/d SRegister_10$1_4/q
+ VSSd VSSd VSSd VSSd VDDd VSSd VSSd VSSd VSSd VSSd out[6] out[4] out[10] out[7] out[5]
+ out[8] qw_NOLclk_0/PHI_2 SRegister_10$1_4/en VDDd qw_NOLclk_0/PHI_1 VSSd SRegister_10$1
XSCHMITT_0 VDDd VSSd SCHMITT_0/IN SCHMITT_0/OUT SCHMITT
.ends

