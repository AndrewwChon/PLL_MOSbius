* Extracted by KLayout with GF180MCU LVS runset on : 13/08/2025 05:13

.SUBCKT asc_9_bit_counter_20250809 vss done vdd a rst d1 d2 d3 d4 d5 d6 d7 d8 d9
M$1 vdd \$56 \$1 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$2 \$1 \$54 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$3 vdd \$52 \$2 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$4 \$2 \$50 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$5 \$3 \$2 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U PD=10.82U
M$7 \$3 \$1 \$4 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U PD=10.82U
M$9 vdd \$4 \$5 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$10 \$5 \$12 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$11 \$6 \$5 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$12 \$105 \$104 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$13 \$216 \$105 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$15 \$217 \$104 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$17 \$217 \$107 \$42 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$19 \$216 \$108 \$42 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$21 vdd \$107 \$108 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$22 \$110 \$109 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$23 \$218 \$110 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$25 \$219 \$109 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$27 \$219 \$112 \$44 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$29 \$218 \$113 \$44 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$31 vdd \$112 \$113 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$32 \$115 \$114 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$33 \$220 \$115 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$35 \$221 \$114 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$37 \$221 \$117 \$46 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$39 \$220 \$118 \$46 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$41 vdd \$117 \$118 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$42 \$120 \$119 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$43 \$222 \$120 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$45 \$223 \$119 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$47 \$223 \$122 \$48 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$49 \$222 \$123 \$48 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$51 vdd \$122 \$123 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$52 \$125 \$124 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$53 \$224 \$125 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$55 \$225 \$124 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$57 \$225 \$127 \$50 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$59 \$224 \$128 \$50 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$61 vdd \$127 \$128 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$62 \$130 \$129 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$63 \$226 \$130 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$65 \$227 \$129 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$67 \$227 \$132 \$52 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$69 \$226 \$133 \$52 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$71 vdd \$132 \$133 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$72 \$135 \$134 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$73 \$228 \$135 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$75 \$229 \$134 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$77 \$229 \$137 \$54 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$79 \$228 \$138 \$54 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$81 vdd \$137 \$138 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$82 \$140 \$139 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$83 \$230 \$140 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$85 \$231 \$139 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$87 \$231 \$142 \$56 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$89 \$230 \$143 \$56 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$91 vdd \$142 \$143 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$92 \$145 \$144 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$93 \$232 \$145 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$95 \$233 \$144 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$97 \$233 \$147 \$58 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$99 \$232 \$148 \$58 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$101 vdd \$147 \$148 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$102 vdd \$48 \$41 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$103 \$41 \$46 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$104 vdd \$44 \$149 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$105 \$149 \$42 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$106 \$234 \$149 vdd vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$108 \$234 \$41 \$12 vdd pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$110 vdd \$58 \$150 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$111 \$150 \$6 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$112 done \$150 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$113 \$758 \$444 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$114 \$444 a vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$115 \$774 \$459 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$116 \$340 \$444 \$339 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$117 vdd \$457 \$340 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$118 \$339 \$758 \$774 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$119 \$457 \$339 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$120 \$340 \$445 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$121 \$341 \$444 \$457 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$122 vdd rst \$445 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$123 vdd \$341 \$459 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$124 \$342 \$758 \$341 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$125 vdd \$459 \$342 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$126 \$459 \$445 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$127 \$107 \$459 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$128 \$104 d1 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$129 \$760 \$446 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$130 \$446 \$107 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$131 \$776 \$461 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$132 \$344 \$446 \$343 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$133 \$343 \$760 \$776 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$134 vdd \$460 \$344 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$135 \$460 \$343 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$136 \$344 \$345 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$137 \$346 \$446 \$460 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$138 vdd rst \$345 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$139 vdd \$346 \$461 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$140 \$347 \$760 \$346 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$141 vdd \$461 \$347 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$142 \$461 \$345 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$143 \$109 d2 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$144 \$112 \$461 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$145 \$762 \$447 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$146 \$447 \$112 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$147 \$778 \$463 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$148 \$349 \$447 \$348 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$149 vdd \$462 \$349 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$150 \$348 \$762 \$778 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$151 \$462 \$348 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$152 \$349 \$350 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$153 \$351 \$447 \$462 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$154 vdd rst \$350 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$155 vdd \$351 \$463 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$156 \$352 \$762 \$351 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$157 vdd \$463 \$352 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$158 \$463 \$350 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$159 \$114 d3 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$160 \$117 \$463 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$161 \$764 \$448 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$162 \$448 \$117 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$163 \$780 \$465 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$164 \$354 \$448 \$353 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$165 \$353 \$764 \$780 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$166 vdd \$464 \$354 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$167 \$464 \$353 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$168 \$354 \$449 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$169 \$355 \$448 \$464 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$170 vdd rst \$449 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$171 vdd \$355 \$465 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$172 \$356 \$764 \$355 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$173 vdd \$465 \$356 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$174 \$465 \$449 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$175 \$119 d4 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$176 \$122 \$465 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$177 \$766 \$450 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$178 \$450 \$122 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$179 \$782 \$467 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$180 \$358 \$450 \$357 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$181 \$357 \$766 \$782 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$182 vdd \$466 \$358 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$183 \$466 \$357 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$184 \$358 \$359 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$185 \$360 \$450 \$466 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$186 vdd rst \$359 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$187 vdd \$360 \$467 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$188 \$361 \$766 \$360 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$189 vdd \$467 \$361 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$190 \$467 \$359 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$191 \$127 \$467 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$192 \$124 d5 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$193 \$768 \$451 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$194 \$451 \$127 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$195 \$784 \$469 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$196 \$363 \$451 \$362 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$197 \$362 \$768 \$784 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$198 vdd \$468 \$363 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$199 \$468 \$362 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$200 \$363 \$364 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$201 \$365 \$451 \$468 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$202 vdd rst \$364 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$203 vdd \$365 \$469 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$204 \$366 \$768 \$365 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$205 vdd \$469 \$366 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$206 \$469 \$364 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$207 \$132 \$469 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$208 \$129 d6 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$209 \$630 \$452 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$210 \$452 \$132 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$211 \$786 \$471 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$212 \$368 \$452 \$367 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$213 \$367 \$630 \$786 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$214 vdd \$470 \$368 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$215 \$470 \$367 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$216 \$368 \$453 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$217 \$369 \$452 \$470 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$218 vdd rst \$453 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$219 vdd \$369 \$471 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$220 \$370 \$630 \$369 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$221 vdd \$471 \$370 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$222 \$471 \$453 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$223 \$134 d7 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$224 \$137 \$471 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$225 \$631 \$454 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$226 \$454 \$137 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$227 \$788 \$473 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$228 \$372 \$454 \$371 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$229 \$371 \$631 \$788 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$230 vdd \$472 \$372 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$231 \$472 \$371 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$232 \$372 \$373 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$233 \$374 \$454 \$472 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$234 vdd rst \$373 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$235 vdd \$374 \$473 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$236 \$375 \$631 \$374 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$237 vdd \$473 \$375 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$238 \$473 \$373 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$239 \$142 \$473 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$240 \$139 d8 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$241 \$772 \$455 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$242 \$455 \$142 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$243 \$790 \$475 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$244 \$377 \$455 \$376 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$245 \$376 \$772 \$790 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$246 vdd \$474 \$377 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$247 \$474 \$376 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$248 \$377 \$378 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$249 \$379 \$455 \$474 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$250 vdd rst \$378 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$251 vdd \$379 \$475 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$252 \$380 \$772 \$379 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$253 vdd \$475 \$380 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$254 \$475 \$378 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$255 \$147 \$475 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$256 \$144 d9 vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$257 \$24 \$56 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$259 \$24 \$54 \$1 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$261 \$25 \$52 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$263 \$25 \$50 \$2 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$265 vss \$2 \$4 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$266 \$4 \$1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$267 \$26 \$4 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U PD=4.74U
M$269 \$26 \$12 \$5 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$271 \$6 \$5 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$272 \$105 \$104 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$273 \$43 \$105 \$42 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$275 \$106 \$104 \$42 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$277 \$43 \$107 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$279 \$106 \$108 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$281 vss \$107 \$108 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$282 \$110 \$109 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$283 \$45 \$110 \$44 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$285 \$111 \$109 \$44 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$287 \$45 \$112 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$289 \$111 \$113 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$291 vss \$112 \$113 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$292 \$115 \$114 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$293 \$47 \$115 \$46 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$295 \$116 \$114 \$46 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$297 \$47 \$117 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$299 \$116 \$118 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$301 vss \$117 \$118 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$302 \$120 \$119 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$303 \$49 \$120 \$48 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$305 \$121 \$119 \$48 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$307 \$49 \$122 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$309 \$121 \$123 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$311 vss \$122 \$123 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$312 \$125 \$124 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$313 \$51 \$125 \$50 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$315 \$126 \$124 \$50 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$317 \$51 \$127 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$319 \$126 \$128 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$321 vss \$127 \$128 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$322 \$130 \$129 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$323 \$53 \$130 \$52 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$325 \$131 \$129 \$52 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$327 \$53 \$132 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$329 \$131 \$133 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$331 vss \$132 \$133 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$332 \$135 \$134 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$333 \$55 \$135 \$54 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$335 \$136 \$134 \$54 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$337 \$55 \$137 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$339 \$136 \$138 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$341 vss \$137 \$138 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$342 \$140 \$139 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$343 \$57 \$140 \$56 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$345 \$141 \$139 \$56 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$347 \$57 \$142 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$349 \$141 \$143 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$351 vss \$142 \$143 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$352 \$145 \$144 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$353 \$59 \$145 \$58 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$355 \$146 \$144 \$58 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$357 \$59 \$147 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$359 \$146 \$148 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$361 vss \$147 \$148 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$362 \$60 \$48 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$364 \$60 \$46 \$41 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$366 \$61 \$44 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$368 \$61 \$42 \$149 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$370 vss \$149 \$12 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$371 \$12 \$41 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$372 \$62 \$58 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$374 \$62 \$6 \$150 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$376 done \$150 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$377 \$758 \$444 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$378 \$444 a vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$379 \$774 \$459 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$380 \$340 \$758 \$339 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$381 \$339 \$444 \$774 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$382 \$549 \$457 \$340 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$384 \$457 \$339 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$385 \$549 \$445 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$387 \$341 \$758 \$457 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$388 vss rst \$445 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$389 \$759 \$341 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$391 \$342 \$444 \$341 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$392 \$759 \$445 \$459 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$394 vss \$459 \$342 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$395 \$107 \$459 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$396 \$104 d1 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$397 \$760 \$446 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$398 \$446 \$107 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$399 \$776 \$461 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$400 \$344 \$760 \$343 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$401 \$550 \$460 \$344 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$403 \$343 \$446 \$776 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$404 \$460 \$343 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$405 \$550 \$345 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$407 \$346 \$760 \$460 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$408 vss rst \$345 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$409 \$761 \$346 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$411 \$347 \$446 \$346 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$412 \$761 \$345 \$461 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$414 vss \$461 \$347 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$415 \$112 \$461 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$416 \$109 d2 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$417 \$762 \$447 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$418 \$447 \$112 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$419 \$778 \$463 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$420 \$349 \$762 \$348 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$421 \$348 \$447 \$778 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$422 \$551 \$462 \$349 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$424 \$462 \$348 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$425 \$551 \$350 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$427 \$351 \$762 \$462 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$428 vss rst \$350 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$429 \$763 \$351 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$431 \$352 \$447 \$351 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$432 \$763 \$350 \$463 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$434 vss \$463 \$352 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$435 \$114 d3 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$436 \$117 \$463 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$437 \$764 \$448 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$438 \$448 \$117 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$439 \$780 \$465 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$440 \$354 \$764 \$353 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$441 \$552 \$464 \$354 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$443 \$353 \$448 \$780 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$444 \$464 \$353 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$445 \$552 \$449 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$447 \$355 \$764 \$464 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$448 vss rst \$449 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$449 \$765 \$355 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$451 \$356 \$448 \$355 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$452 \$765 \$449 \$465 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$454 vss \$465 \$356 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$455 \$122 \$465 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$456 \$119 d4 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$457 \$766 \$450 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$458 \$450 \$122 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$459 \$782 \$467 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$460 \$358 \$766 \$357 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$461 \$357 \$450 \$782 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$462 \$553 \$466 \$358 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$464 \$466 \$357 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$465 \$553 \$359 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$467 \$360 \$766 \$466 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$468 vss rst \$359 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$469 \$767 \$360 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$471 \$361 \$450 \$360 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$472 \$767 \$359 \$467 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$474 vss \$467 \$361 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$475 \$127 \$467 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$476 \$124 d5 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$477 \$768 \$451 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$478 \$451 \$127 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$479 \$784 \$469 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$480 \$363 \$768 \$362 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$481 \$362 \$451 \$784 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$482 \$554 \$468 \$363 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$484 \$468 \$362 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$485 \$554 \$364 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$487 \$365 \$768 \$468 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$488 vss rst \$364 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$489 \$769 \$365 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$491 \$366 \$451 \$365 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$492 \$769 \$364 \$469 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$494 vss \$469 \$366 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$495 \$129 d6 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$496 \$132 \$469 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$497 \$630 \$452 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$498 \$452 \$132 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$499 \$786 \$471 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$500 \$368 \$630 \$367 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$501 \$367 \$452 \$786 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$502 \$555 \$470 \$368 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$504 \$470 \$367 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$505 \$555 \$453 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$507 \$369 \$630 \$470 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$508 vss rst \$453 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$509 \$770 \$369 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$511 \$370 \$452 \$369 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$512 \$770 \$453 \$471 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$514 vss \$471 \$370 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$515 \$137 \$471 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$516 \$134 d7 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$517 \$631 \$454 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$518 \$454 \$137 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$519 \$788 \$473 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$520 \$372 \$631 \$371 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$521 \$371 \$454 \$788 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$522 \$556 \$472 \$372 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$524 \$472 \$371 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$525 \$556 \$373 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$527 \$374 \$631 \$472 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$528 vss rst \$373 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$529 \$771 \$374 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$531 \$375 \$454 \$374 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$532 \$771 \$373 \$473 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$534 vss \$473 \$375 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$535 \$142 \$473 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$536 \$139 d8 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$537 \$772 \$455 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$538 \$455 \$142 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$539 \$790 \$475 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$540 \$377 \$772 \$376 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$541 \$557 \$474 \$377 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$543 \$376 \$455 \$790 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$544 \$474 \$376 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$545 \$557 \$378 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$547 \$379 \$772 \$474 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$548 vss rst \$378 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$549 \$773 \$379 vss vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$551 \$380 \$455 \$379 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$552 \$773 \$378 \$475 vss nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U
+ PD=4.74U
M$554 vss \$475 \$380 vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$555 \$147 \$475 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$556 \$144 d9 vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
.ENDS asc_9_bit_counter_20250809
