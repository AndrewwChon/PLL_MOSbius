* Extracted by KLayout with GF180MCU LVS runset on : 02/08/2025 04:57

.SUBCKT asc_dff_rst vdd clkn|clkp|out ins clkn|clkp|in|out in|ind|ins A|B|out
+ B|ind|ins ins|out A|ind|out clk|in in|rst Qb|in vss Q|out D
M$1 vdd A|ind|out ins vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$2 ins A|B|out vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$3 clkn|clkp|in|out clk|in vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$4 clkn|clkp|out clkn|clkp|in|out vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$5 vdd in|rst A|B|out vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$6 vdd Qb|in ins|out vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$7 ins clkn|clkp|in|out in|ind|ins vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$8 ins|out clkn|clkp|out B|ind|ins vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$9 in|ind|ins clkn|clkp|out \$49 vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$10 B|ind|ins clkn|clkp|in|out A|ind|out vdd pfet_03v3 L=0.5U W=3U AS=1.95P
+ AD=1.95P PS=7.3U PD=7.3U
M$11 \$49 D vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$12 A|ind|out in|ind|ins vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P
+ PS=7.3U PD=7.3U
M$13 Q|out Qb|in vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$14 vdd B|ind|ins Qb|in vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$15 Qb|in A|B|out vdd vdd pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U
+ PD=7.3U
M$16 ins clkn|clkp|out in|ind|ins vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$17 ins|out clkn|clkp|in|out B|ind|ins vss nfet_03v3 L=0.5U W=1U AS=0.61P
+ AD=0.61P PS=3.22U PD=3.22U
M$18 clkn|clkp|in|out clk|in vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$19 clkn|clkp|out clkn|clkp|in|out vss vss nfet_03v3 L=0.5U W=1U AS=0.61P
+ AD=0.61P PS=3.22U PD=3.22U
M$20 vss in|rst A|B|out vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$21 vss Qb|in ins|out vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$22 \$32 A|ind|out ins vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$23 vss A|B|out \$32 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$24 \$48 B|ind|ins vss vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$25 Qb|in A|B|out \$48 vss nfet_03v3 L=0.5U W=2U AS=1.22P AD=1.22P PS=5.22U
+ PD=5.22U
M$26 \$49 D vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$27 A|ind|out in|ind|ins vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P
+ PS=3.22U PD=3.22U
M$28 Q|out Qb|in vss vss nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U
+ PD=3.22U
M$29 in|ind|ins clkn|clkp|in|out \$49 vss nfet_03v3 L=0.5U W=1U AS=0.61P
+ AD=0.61P PS=3.22U PD=3.22U
M$30 B|ind|ins clkn|clkp|out A|ind|out vss nfet_03v3 L=0.5U W=1U AS=0.61P
+ AD=0.61P PS=3.22U PD=3.22U
.ENDS asc_dff_rst
