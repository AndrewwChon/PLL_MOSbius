* Extracted by KLayout with GF180MCU LVS runset on : 09/08/2025 20:59

.SUBCKT asc_XNOR VSS OUT A B VDD
M$1 \$9 A VDD VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$2 \$20 \$9 VDD VDD pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U PD=10.82U
M$4 \$21 A VDD VDD pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U PD=10.82U
M$6 \$21 B OUT VDD pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U PD=10.82U
M$8 \$20 \$12 OUT VDD pfet_03v3 L=0.5U W=6U AS=2.73P AD=2.73P PS=10.82U
+ PD=10.82U
M$10 VDD B \$12 VDD pfet_03v3 L=0.5U W=3U AS=1.95P AD=1.95P PS=7.3U PD=7.3U
M$11 \$9 A VSS VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
M$12 \$3 \$9 OUT VSS nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U PD=4.74U
M$14 \$10 A OUT VSS nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U PD=4.74U
M$16 \$3 B VSS VSS nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U PD=4.74U
M$18 \$10 \$12 VSS VSS nfet_03v3 L=0.5U W=2U AS=0.87P AD=0.87P PS=4.74U PD=4.74U
M$20 VSS B \$12 VSS nfet_03v3 L=0.5U W=1U AS=0.61P AD=0.61P PS=3.22U PD=3.22U
.ENDS asc_XNOR
