** sch_path: /foss/designs/libs/qw_core_analog/PCP1248Xflatten/PCP1248Xflatten.sch
.subckt PCP1248Xflatten vdd vss vin iref200u out up down s0 s1 s2 s3
*.PININFO vdd:B vss:B vin:B iref200u:B out:B up:B down:B s0:B s1:B s2:B s3:B
M25 net1 s0b vss vss nfet_03v3 L=0.28u W=2u nf=1 m=1
M26 net2 net1 vss vss nfet_03v3 L=0.5u W=8u nf=4 m=1
M27 net14 vb1 net2 vss nfet_03v3 L=0.5u W=8u nf=4 m=1
M28 net3 s1b vss vss nfet_03v3 L=0.28u W=2u nf=1 m=1
M29 net4 net3 vss vss nfet_03v3 L=0.5u W=8u nf=4 m=2
M30 net14 vb1 net4 vss nfet_03v3 L=0.5u W=8u nf=4 m=2
M31 net5 s2b vss vss nfet_03v3 L=0.28u W=2u nf=1 m=1
M32 net6 net5 vss vss nfet_03v3 L=0.5u W=8u nf=4 m=4
M33 net14 vb1 net6 vss nfet_03v3 L=0.5u W=8u nf=4 m=4
M34 net13 vb2 net7 vdd pfet_03v3 L=0.5u W=20u nf=8 m=1
M35 net7 net8 vdd vdd pfet_03v3 L=0.5u W=20u nf=8 m=1
M36 net8 s0 vdd vdd pfet_03v3 L=0.28u W=2u nf=1 m=1
M37 net13 vb2 net9 vdd pfet_03v3 L=0.5u W=20u nf=8 m=2
M38 net9 net10 vdd vdd pfet_03v3 L=0.5u W=20u nf=8 m=2
M39 net10 s1 vdd vdd pfet_03v3 L=0.28u W=2u nf=1 m=1
M40 net13 vb2 net11 vdd pfet_03v3 L=0.5u W=20u nf=8 m=4
M41 net11 net12 vdd vdd pfet_03v3 L=0.5u W=20u nf=8 m=4
M42 net12 s2 vdd vdd pfet_03v3 L=0.28u W=2u nf=1 m=1
M43 out down net14 vss nfet_03v3 L=0.28u W=8u nf=1 m=1
M44 out up net13 vdd pfet_03v3 L=0.28u W=20u nf=1 m=1
M15 net16 gatep vdd vdd pfet_03v3 L=0.5u W=20u nf=8 m=1
M16 gatep vb2 net16 vdd pfet_03v3 L=0.5u W=20u nf=8 m=1
M23 net15 gaten vss vss nfet_03v3 L=0.5u W=8u nf=4 m=1
M24 gatep vb1 net15 vss nfet_03v3 L=0.5u W=8u nf=4 m=1
M45 vb2 gaten vss vss nfet_03v3 L=0.5u W=4u nf=4 m=2
M46 vb2 vb2 vdd vdd pfet_03v3 L=0.5u W=2.5u nf=2 m=2
M47 vb1 vb2 vdd vdd pfet_03v3 L=0.5u W=2.5u nf=2 m=2
M48 vb1 vb1 vss vss nfet_03v3 L=0.5u W=2u nf=2 m=1
M49 net17 gaten vss vss nfet_03v3 L=0.5u W=4u nf=4 m=2
M50 vdd vb1 net17 vss nfet_03v3 L=0.5u W=8u nf=1 m=1
x8 vdd iref200u vdd vin gaten vss OTAforChargePump
x9 s0 vdd s0b vss inv1u05u
x10 s1 vdd s1b vss inv1u05u
x11 s2 vdd s2b vss inv1u05u
M1 net18 s3b vss vss nfet_03v3 L=0.28u W=2u nf=1 m=1
M2 net19 net18 vss vss nfet_03v3 L=0.5u W=8u nf=4 m=8
M3 net14 vb1 net19 vss nfet_03v3 L=0.5u W=8u nf=4 m=8
M4 net13 vb2 net20 vdd pfet_03v3 L=0.5u W=20u nf=8 m=8
M5 net20 net21 vdd vdd pfet_03v3 L=0.5u W=20u nf=8 m=8
M6 net21 s3 vdd vdd pfet_03v3 L=0.28u W=2u nf=1 m=1
x13 s3 vdd s3b vss inv1u05u
M7 vss vss vss vss nfet_03v3 L=0.5u W=2u nf=2 m=2
M8 vdd vdd vdd vdd pfet_03v3 L=0.5u W=2.5u nf=2 m=2
M9 vdd vdd vdd vdd pfet_03v3 L=0.5u W=10u nf=4 m=6
M10 vdd vdd vdd vdd pfet_03v3 L=0.5u W=20u nf=8 m=2
M11 net13 net13 net13 vdd pfet_03v3 L=0.5u W=10u nf=4 m=5
M12 net13 net13 net13 vdd pfet_03v3 L=0.5u W=20u nf=8 m=2
M13 gatep gatep gatep vdd pfet_03v3 L=0.5u W=10u nf=4 m=1
M14 vss vss vss vss nfet_03v3 L=0.5u W=4u nf=2 m=6
M17 vss vss vss vss nfet_03v3 L=0.5u W=8u nf=4 m=2
M18 net14 net14 net14 vss nfet_03v3 L=0.5u W=4u nf=2 m=5
M19 net14 net14 net14 vss nfet_03v3 L=0.5u W=8u nf=4 m=2
M20 gatep gatep gatep vss nfet_03v3 L=0.5u W=4u nf=2 m=1
x14 vdd s0b gaten net1 vss s0 TG
x1 vdd s1b gaten net3 vss s1 TG
x2 vdd s2b gaten net5 vss s2 TG
x3 vdd s3b gaten net18 vss s3 TG
x4 vdd s0b gatep net8 vss s0 TG
x5 vdd s1b gatep net10 vss s1 TG
x6 vdd s2b gatep net12 vss s2 TG
x7 vdd s3b gatep net21 vss s3 TG
.ends

* expanding   symbol:  libs/qw_core_analog/OTAforChargePump/OTAforChargePump.sym # of pins=6
** sym_path: /foss/designs/libs/qw_core_analog/OTAforChargePump/OTAforChargePump.sym
** sch_path: /foss/designs/libs/qw_core_analog/OTAforChargePump/OTAforChargePump.sch
.subckt OTAforChargePump vdd iref inp inn out vss
*.PININFO inp:B inn:B vdd:B vss:B out:B iref:B
M8 iref iref vdd vdd pfet_03v3 L=0.28u W=10u nf=4 m=4
M1 net1 iref vdd vdd pfet_03v3 L=0.28u W=10u nf=4 m=4
M2 net2 inp net1 vdd pfet_03v3 L=0.28u W=10u nf=4 m=2
M3 out inn net1 vdd pfet_03v3 L=0.28u W=10u nf=4 m=2
M4 net2 net2 vss vss nfet_03v3 L=0.28u W=4u nf=2 m=2
M5 out net2 vss vss nfet_03v3 L=0.28u W=4u nf=2 m=2
M6 vdd vdd vdd vdd pfet_03v3 L=0.28u W=5u nf=2 m=4
M7 vss vss vss vss nfet_03v3 L=0.28u W=8u nf=4 m=2
M9 net1 net1 net1 vdd pfet_03v3 L=0.28u W=5u nf=2 m=2
.ends


* expanding   symbol:  libs/xp_core_analog/inv1u05u/inv1u05u.sym # of pins=4
** sym_path: /foss/designs/libs/xp_core_analog/inv1u05u/inv1u05u.sym
** sch_path: /foss/designs/libs/xp_core_analog/inv1u05u/inv1u05u.sch
.subckt inv1u05u in vdd out vss
*.PININFO in:B out:B vss:B vdd:B
M1 out in vdd vdd pfet_03v3 L=0.5u W=3.0u nf=1 m=1
M2 out in vss vss nfet_03v3 L=0.5u W=1.0u nf=1 m=1
.ends


* expanding   symbol:  libs/qw_core_analog/TG/TG.sym # of pins=6
** sym_path: /foss/designs/libs/qw_core_analog/TG/TG.sym
** sch_path: /foss/designs/libs/qw_core_analog/TG/TG.sch
.subckt TG vdd clkp ind ins vss clkn
*.PININFO ind:B ins:B clkn:B clkp:B vdd:B vss:B
M1 ind clkp ins vdd pfet_03v3 L=0.28u W=2u nf=1 m=1
M2 ind clkn ins vss nfet_03v3 L=0.28u W=2u nf=1 m=1
.ends

