* Extracted by KLayout with GF180MCU LVS runset on : 29/08/2025 01:57

.SUBCKT SCHMITT VSS IN VDD OUT vss
M$1 VSS OUT \$10 VDD pfet_03v3 L=0.28U W=2U AS=1.3P AD=1.3P PS=5.3U PD=5.3U
M$2 \$10 IN VDD VDD pfet_03v3 L=0.28U W=4U AS=2.6P AD=2.6P PS=9.3U PD=9.3U
M$3 OUT IN \$10 VDD pfet_03v3 L=0.28U W=4U AS=2.6P AD=2.6P PS=9.3U PD=9.3U
M$4 \$3 IN VSS vss nfet_03v3 L=0.28U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$5 OUT IN \$3 vss nfet_03v3 L=0.28U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
M$6 VDD OUT \$3 vss nfet_03v3 L=0.28U W=2U AS=1.22P AD=1.22P PS=5.22U PD=5.22U
.ENDS SCHMITT
