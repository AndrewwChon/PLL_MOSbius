* NGSPICE file created from top_level_20250921.ext - technology: gf180mcuD

.subckt cap_nmos$2 a_88_n92# a_0_0#
X0 a_88_n92# a_0_0# cap_nmos_03v3 c_width=10u c_length=10u
.ends

.subckt DECAP_SC$1 a_n313_2257# vdd vss
Xcap_nmos$2_0 vdd vss cap_nmos$2
Xcap_nmos$2_1 vdd vss cap_nmos$2
Xcap_nmos$2_2 vdd vss cap_nmos$2
Xcap_nmos$2_3 vdd vss cap_nmos$2
.ends

.subckt DECAP_LARGE vdd vss
XDECAP_SC$1_121 vss vdd vss DECAP_SC$1
XDECAP_SC$1_110 vss vdd vss DECAP_SC$1
XDECAP_SC$1_70 vss vdd vss DECAP_SC$1
XDECAP_SC$1_81 vss vdd vss DECAP_SC$1
XDECAP_SC$1_92 vss vdd vss DECAP_SC$1
XDECAP_SC$1_122 vss vdd vss DECAP_SC$1
XDECAP_SC$1_100 vss vdd vss DECAP_SC$1
XDECAP_SC$1_111 vss vdd vss DECAP_SC$1
XDECAP_SC$1_71 vss vdd vss DECAP_SC$1
XDECAP_SC$1_60 vss vdd vss DECAP_SC$1
XDECAP_SC$1_93 vss vdd vss DECAP_SC$1
XDECAP_SC$1_82 vss vdd vss DECAP_SC$1
XDECAP_SC$1_123 vss vdd vss DECAP_SC$1
XDECAP_SC$1_101 vss vdd vss DECAP_SC$1
XDECAP_SC$1_112 DECAP_SC$1_112/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_50 vss vdd vss DECAP_SC$1
XDECAP_SC$1_72 DECAP_SC$1_72/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_94 vss vdd vss DECAP_SC$1
XDECAP_SC$1_61 vss vdd vss DECAP_SC$1
XDECAP_SC$1_83 vss vdd vss DECAP_SC$1
XDECAP_SC$1_102 DECAP_SC$1_102/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_124 vss vdd vss DECAP_SC$1
XDECAP_SC$1_113 vss vdd vss DECAP_SC$1
XDECAP_SC$1_40 DECAP_SC$1_40/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_51 vss vdd vss DECAP_SC$1
XDECAP_SC$1_73 vss vdd vss DECAP_SC$1
XDECAP_SC$1_95 vss vdd vss DECAP_SC$1
XDECAP_SC$1_62 vss vdd vss DECAP_SC$1
XDECAP_SC$1_84 vss vdd vss DECAP_SC$1
XDECAP_SC$1_103 DECAP_SC$1_103/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_125 vss vdd vss DECAP_SC$1
XDECAP_SC$1_114 vss vdd vss DECAP_SC$1
XDECAP_SC$1_52 DECAP_SC$1_52/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_41 DECAP_SC$1_41/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_30 vss vdd vss DECAP_SC$1
XDECAP_SC$1_96 DECAP_SC$1_96/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_63 vss vdd vss DECAP_SC$1
XDECAP_SC$1_74 vss vdd vss DECAP_SC$1
XDECAP_SC$1_85 vss vdd vss DECAP_SC$1
XDECAP_SC$1_104 DECAP_SC$1_104/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_115 vss vdd vss DECAP_SC$1
XDECAP_SC$1_64 vss vdd vss DECAP_SC$1
XDECAP_SC$1_42 vss vdd vss DECAP_SC$1
XDECAP_SC$1_31 vss vdd vss DECAP_SC$1
XDECAP_SC$1_20 vss vdd vss DECAP_SC$1
XDECAP_SC$1_97 vss vdd vss DECAP_SC$1
XDECAP_SC$1_53 vss vdd vss DECAP_SC$1
XDECAP_SC$1_75 vss vdd vss DECAP_SC$1
XDECAP_SC$1_86 vss vdd vss DECAP_SC$1
XDECAP_SC$1_105 DECAP_SC$1_105/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_116 vss vdd vss DECAP_SC$1
XDECAP_SC$1_65 vss vdd vss DECAP_SC$1
XDECAP_SC$1_43 vss vdd vss DECAP_SC$1
XDECAP_SC$1_54 vss vdd vss DECAP_SC$1
XDECAP_SC$1_21 vss vdd vss DECAP_SC$1
XDECAP_SC$1_10 vss vdd vss DECAP_SC$1
XDECAP_SC$1_98 vss vdd vss DECAP_SC$1
XDECAP_SC$1_32 DECAP_SC$1_32/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_76 vss vdd vss DECAP_SC$1
XDECAP_SC$1_87 vss vdd vss DECAP_SC$1
XDECAP_SC$1_106 DECAP_SC$1_106/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_117 vss vdd vss DECAP_SC$1
XDECAP_SC$1_66 vss vdd vss DECAP_SC$1
XDECAP_SC$1_44 DECAP_SC$1_44/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_88 vss vdd vss DECAP_SC$1
XDECAP_SC$1_55 vss vdd vss DECAP_SC$1
XDECAP_SC$1_22 vss vdd vss DECAP_SC$1
XDECAP_SC$1_11 vss vdd vss DECAP_SC$1
XDECAP_SC$1_99 vss vdd vss DECAP_SC$1
XDECAP_SC$1_33 vss vdd vss DECAP_SC$1
XDECAP_SC$1_77 vss vdd vss DECAP_SC$1
XDECAP_SC$1_107 DECAP_SC$1_107/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_118 vss vdd vss DECAP_SC$1
XDECAP_SC$1_67 vss vdd vss DECAP_SC$1
XDECAP_SC$1_89 vss vdd vss DECAP_SC$1
XDECAP_SC$1_56 vss vdd vss DECAP_SC$1
XDECAP_SC$1_23 vss vdd vss DECAP_SC$1
XDECAP_SC$1_12 DECAP_SC$1_12/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_34 vss vdd vss DECAP_SC$1
XDECAP_SC$1_45 DECAP_SC$1_45/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_78 vss vdd vss DECAP_SC$1
XDECAP_SC$1_108 DECAP_SC$1_108/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_119 vss vdd vss DECAP_SC$1
XDECAP_SC$1_46 vss vdd vss DECAP_SC$1
XDECAP_SC$1_68 vss vdd vss DECAP_SC$1
XDECAP_SC$1_57 vss vdd vss DECAP_SC$1
XDECAP_SC$1_24 vss vdd vss DECAP_SC$1
XDECAP_SC$1_13 vss vdd vss DECAP_SC$1
XDECAP_SC$1_35 vss vdd vss DECAP_SC$1
XDECAP_SC$1_79 vss vdd vss DECAP_SC$1
XDECAP_SC$1_109 DECAP_SC$1_109/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_47 vss vdd vss DECAP_SC$1
XDECAP_SC$1_69 vss vdd vss DECAP_SC$1
XDECAP_SC$1_25 vss vdd vss DECAP_SC$1
XDECAP_SC$1_14 vss vdd vss DECAP_SC$1
XDECAP_SC$1_58 vss vdd vss DECAP_SC$1
XDECAP_SC$1_36 vss vdd vss DECAP_SC$1
XDECAP_SC$1_48 vss vdd vss DECAP_SC$1
XDECAP_SC$1_26 vss vdd vss DECAP_SC$1
XDECAP_SC$1_15 vss vdd vss DECAP_SC$1
XDECAP_SC$1_59 DECAP_SC$1_59/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_37 vss vdd vss DECAP_SC$1
XDECAP_SC$1_49 vss vdd vss DECAP_SC$1
XDECAP_SC$1_0 vss vdd vss DECAP_SC$1
XDECAP_SC$1_27 vss vdd vss DECAP_SC$1
XDECAP_SC$1_16 vss vdd vss DECAP_SC$1
XDECAP_SC$1_38 vss vdd vss DECAP_SC$1
XDECAP_SC$1_1 vss vdd vss DECAP_SC$1
XDECAP_SC$1_28 vss vdd vss DECAP_SC$1
XDECAP_SC$1_17 vss vdd vss DECAP_SC$1
XDECAP_SC$1_39 vss vdd vss DECAP_SC$1
XDECAP_SC$1_2 DECAP_SC$1_2/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_29 vss vdd vss DECAP_SC$1
XDECAP_SC$1_18 vss vdd vss DECAP_SC$1
XDECAP_SC$1_3 DECAP_SC$1_3/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_19 vss vdd vss DECAP_SC$1
XDECAP_SC$1_4 DECAP_SC$1_4/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_5 DECAP_SC$1_5/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_6 DECAP_SC$1_6/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_7 DECAP_SC$1_7/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_8 DECAP_SC$1_8/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_9 DECAP_SC$1_9/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_90 DECAP_SC$1_90/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_120 DECAP_SC$1_120/a_n313_2257# vdd vss DECAP_SC$1
XDECAP_SC$1_80 vss vdd vss DECAP_SC$1
XDECAP_SC$1_91 DECAP_SC$1_91/a_n313_2257# vdd vss DECAP_SC$1
.ends

.subckt ppolyf_u_resistor$9 a_n376_0# a_5400_0# a_n132_0#
X0 a_n132_0# a_5400_0# a_n376_0# ppolyf_u r_width=1u r_length=27u
.ends

.subckt ppolyf_u_resistor$8 a_n376_0# a_1100_0# a_n132_0#
X0 a_n132_0# a_1100_0# a_n376_0# ppolyf_u r_width=40u r_length=5.5u
.ends

.subckt diode_pd2nw$1 w_n224_n86# a_0_0#
D0 a_0_0# w_n224_n86# diode_pd2nw_03v3 pj=40u area=99.99999p
.ends

.subckt diode_nd2ps$1 a_n168_0# a_0_0#
D0 a_n168_0# a_0_0# diode_nd2ps_03v3 pj=40u area=99.99999p
.ends

.subckt io_secondary_3p3 ASIG3V3 VDD VSS to_gate
Xppolyf_u_resistor$8_0 VSS ASIG3V3 to_gate ppolyf_u_resistor$8
Xdiode_pd2nw$1_0 VDD to_gate diode_pd2nw$1
Xdiode_pd2nw$1_1 VDD to_gate diode_pd2nw$1
Xdiode_pd2nw$1_3 VDD to_gate diode_pd2nw$1
Xdiode_pd2nw$1_2 VDD to_gate diode_pd2nw$1
Xdiode_nd2ps$1_0 VSS to_gate diode_nd2ps$1
Xdiode_nd2ps$1_1 VSS to_gate diode_nd2ps$1
Xdiode_nd2ps$1_3 VSS to_gate diode_nd2ps$1
Xdiode_nd2ps$1_2 VSS to_gate diode_nd2ps$1
.ends

.subckt ppolyf_u_resistor a_n376_0# a_1100_0# a_n132_0#
X0 a_n132_0# a_1100_0# a_n376_0# ppolyf_u r_width=40u r_length=5.5u
.ends

.subckt nfet$465 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$463 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$461 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$439 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$437 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$435 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$464 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$462 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$438 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$436 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt asc_hysteresis_buffer$9 vss in vdd out
Xnfet$465_0 m1_1156_42# vss m1_884_42# vss nfet$465
Xnfet$463_0 in vss m1_348_648# vss nfet$463
Xnfet$461_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$461
Xpfet$439_0 vdd vdd m1_884_42# m1_1156_42# pfet$439
Xpfet$437_0 vdd vdd m1_348_648# in pfet$437
Xpfet$435_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd
+ m1_884_42# m1_884_42# pfet$435
Xnfet$464_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$464
Xnfet$462_0 m1_348_648# vss m1_884_42# vss nfet$462
Xpfet$438_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$438
Xpfet$436_0 vdd vdd m1_884_42# m1_348_648# pfet$436
.ends

.subckt pfet$440 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=2.6p pd=9.3u as=2.6p ps=9.3u w=4u l=0.28u
.ends

.subckt nfet$466 a_n84_0# a_94_0# a_30_460# VSUBS
X0 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$441 a_28_460# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_460# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt nfet$467 a_30_n132# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt SCHMITT$4 VDD VSS IN OUT
Xpfet$440_0 IN VDD m1_596_1544# OUT pfet$440
Xnfet$466_0 m1_592_402# OUT IN VSS nfet$466
Xpfet$440_1 IN VDD VDD m1_596_1544# pfet$440
Xnfet$466_1 VSS m1_592_402# IN VSS nfet$466
Xpfet$441_0 OUT VDD m1_596_1544# VSS pfet$441
Xnfet$467_0 OUT m1_592_402# VDD VSS nfet$467
.ends

.subckt nfet$470 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$444 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$442 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt nfet$468 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt nfet$471 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$445 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$469 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt pfet$443 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt qw_NOLclk$2 CLK VDDd VSSd PHI_1 PHI_2
Xnfet$470_0 m1_11601_71# VSSd PHI_1 VSSd nfet$470
Xnfet$470_1 m1_11161_409# VSSd m1_11379_n171# VSSd nfet$470
Xnfet$470_2 m1_11601_2380# VSSd PHI_2 VSSd nfet$470
Xnfet$470_3 CLK VSSd m1_11161_409# VSSd nfet$470
Xpfet$444_0 VDDd VDDd PHI_1 m1_11601_71# pfet$444
Xpfet$444_1 VDDd VDDd m1_11379_n171# m1_11161_409# pfet$444
Xpfet$444_2 VDDd VDDd PHI_2 m1_11601_2380# pfet$444
Xpfet$444_3 VDDd VDDd m1_11161_409# CLK pfet$444
Xpfet$442_0 VDDd VDDd m1_13930_233# PHI_1 pfet$442
Xpfet$442_1 VDDd VDDd m1_13930_1818# PHI_2 pfet$442
Xnfet$468_1 PHI_2 VSSd m1_13930_1818# VSSd nfet$468
Xnfet$468_0 PHI_1 VSSd m1_13930_233# VSSd nfet$468
Xnfet$471_0 m1_12351_431# m1_12351_431# m1_11601_71# m1_11601_71# m1_11837_749# VSSd
+ nfet$471
Xnfet$471_1 m1_11379_n171# m1_11379_n171# VSSd VSSd m1_11837_749# VSSd nfet$471
Xnfet$471_2 m1_12351_2064# m1_12351_2064# m1_11601_2380# m1_11601_2380# m1_11837_1708#
+ VSSd nfet$471
Xnfet$471_3 m1_11161_409# m1_11161_409# VSSd VSSd m1_11837_1708# VSSd nfet$471
Xpfet$445_0 VDDd m1_11601_71# VDDd m1_11379_n171# pfet$445
Xpfet$445_1 VDDd VDDd m1_11601_71# m1_12351_431# pfet$445
Xpfet$445_2 VDDd m1_11601_2380# VDDd m1_11161_409# pfet$445
Xpfet$445_3 VDDd VDDd m1_11601_2380# m1_12351_2064# pfet$445
Xnfet$469_0 m1_12351_2064# m1_15103_233# VSSd VSSd nfet$469
Xpfet$443_0 m1_12351_2064# VDDd VDDd m1_15103_233# pfet$443
Xnfet$469_1 m1_15103_233# m1_13930_233# VSSd VSSd nfet$469
Xpfet$443_1 m1_15103_233# VDDd VDDd m1_13930_233# pfet$443
Xpfet$443_2 m1_12351_431# VDDd VDDd m1_15103_1818# pfet$443
Xpfet$443_3 m1_15103_1818# VDDd VDDd m1_13930_1818# pfet$443
Xnfet$469_2 m1_12351_431# m1_15103_1818# VSSd VSSd nfet$469
Xnfet$469_3 m1_15103_1818# m1_13930_1818# VSSd VSSd nfet$469
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__or2_1$4 A1 A2 VDD VSS Z VNW VPW
X0 a_255_756# A1 a_67_756# VNW pfet_05v0 ad=0.2379p pd=1.435u as=0.4026p ps=2.71u w=0.915u l=0.5u
X1 VSS A2 a_67_756# VPW nfet_05v0 ad=0.3828p pd=2.08u as=0.1716p ps=1.18u w=0.66u l=0.6u
X2 VDD A2 a_255_756# VNW pfet_05v0 ad=0.57645p pd=2.69u as=0.2379p ps=1.435u w=0.915u l=0.5u
X3 Z a_67_756# VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.3828p ps=2.08u w=1.32u l=0.6u
X4 Z a_67_756# VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.57645p ps=2.69u w=1.83u l=0.5u
X5 a_67_756# A1 VSS VPW nfet_05v0 ad=0.1716p pd=1.18u as=0.2904p ps=2.2u w=0.66u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1$4 I VDD VSS ZN VNW VPW
X0 ZN I VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__latq_1$5 D E Q VDD VSS VNW VPW
X0 VSS a_1020_652# Q VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X1 a_504_110# a_36_92# VDD VNW pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X2 VDD a_1020_652# Q VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X3 a_1264_107# a_36_92# a_1020_652# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X4 VSS E a_36_92# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X5 VSS a_1364_532# a_1264_107# VPW nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X6 VDD E a_36_92# VNW pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X7 VDD a_1364_532# a_1224_652# VNW pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X8 a_872_652# D VDD VNW pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X9 a_1364_532# a_1020_652# VDD VNW pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X10 a_1020_652# a_504_110# a_872_107# VPW nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X11 a_872_107# D VSS VPW nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X12 a_1020_652# a_36_92# a_872_652# VNW pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X13 a_504_110# a_36_92# VSS VPW nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X14 a_1364_532# a_1020_652# VSS VPW nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X15 a_1224_652# a_504_110# a_1020_652# VNW pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt DFF_2phase_1$4 VDDd PHI_2 PHI_1 D Q VSSd
Xgf180mcu_fd_sc_mcu9t5v0__latq_1$5_0 gf180mcu_fd_sc_mcu9t5v0__latq_1$5_1/Q PHI_2 Q
+ VDDd VSSd VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1$5
Xgf180mcu_fd_sc_mcu9t5v0__latq_1$5_1 D PHI_1 gf180mcu_fd_sc_mcu9t5v0__latq_1$5_1/Q
+ VDDd VSSd VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1$5
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__and2_1$4 A1 A2 VDD VSS Z VNW VPW
X0 VDD A2 a_36_201# VNW pfet_05v0 ad=0.5054p pd=2.57u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1 a_244_201# A1 a_36_201# VPW nfet_05v0 ad=0.1056p pd=0.98u as=0.2904p ps=2.2u w=0.66u l=0.6u
X2 Z a_36_201# VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.3894p ps=2.06u w=1.32u l=0.6u
X3 Z a_36_201# VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.5054p ps=2.57u w=1.83u l=0.5u
X4 VSS A2 a_244_201# VPW nfet_05v0 ad=0.3894p pd=2.06u as=0.1056p ps=0.98u w=0.66u l=0.6u
X5 a_36_201# A1 VDD VNW pfet_05v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.5u
.ends

.subckt Register_unitcell$3 VDDd out q en default d phi2 phi1 VSSd
Xgf180mcu_fd_sc_mcu9t5v0__or2_1$4_0 gf180mcu_fd_sc_mcu9t5v0__or2_1$4_0/A1 gf180mcu_fd_sc_mcu9t5v0__or2_1$4_0/A2
+ VDDd VSSd out VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1$4
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$4_0 en VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1$4_0/ZN
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1$4
XDFF_2phase_1$4_0 VDDd phi2 phi1 d q VSSd DFF_2phase_1$4
Xgf180mcu_fd_sc_mcu9t5v0__and2_1$4_0 gf180mcu_fd_sc_mcu9t5v0__inv_1$4_0/ZN default
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1$4_0/A1 VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1$4
Xgf180mcu_fd_sc_mcu9t5v0__and2_1$4_1 q en VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1$4_0/A2
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1$4
.ends

.subckt SRegister_10$2 out[1] out[2] out[3] out[5] out[8] d default10 default9 default8
+ default7 default6 default5 default4 default3 default2 default1 out[9] out[6] out[4]
+ out[10] en out[7] q phi2 VDDd VSSd phi1
XRegister_unitcell$3_0 VDDd out[2] Register_unitcell$3_7/d en default2 Register_unitcell$3_6/q
+ phi2 phi1 VSSd Register_unitcell$3
XRegister_unitcell$3_1 VDDd out[6] Register_unitcell$3_2/d en default6 Register_unitcell$3_9/q
+ phi2 phi1 VSSd Register_unitcell$3
XRegister_unitcell$3_2 VDDd out[7] Register_unitcell$3_3/d en default7 Register_unitcell$3_2/d
+ phi2 phi1 VSSd Register_unitcell$3
XRegister_unitcell$3_3 VDDd out[8] Register_unitcell$3_4/d en default8 Register_unitcell$3_3/d
+ phi2 phi1 VSSd Register_unitcell$3
XRegister_unitcell$3_4 VDDd out[9] Register_unitcell$3_5/d en default9 Register_unitcell$3_4/d
+ phi2 phi1 VSSd Register_unitcell$3
XRegister_unitcell$3_5 VDDd out[10] q en default10 Register_unitcell$3_5/d phi2 phi1
+ VSSd Register_unitcell$3
XRegister_unitcell$3_6 VDDd out[1] Register_unitcell$3_6/q en default1 d phi2 phi1
+ VSSd Register_unitcell$3
XRegister_unitcell$3_7 VDDd out[3] Register_unitcell$3_8/d en default3 Register_unitcell$3_7/d
+ phi2 phi1 VSSd Register_unitcell$3
XRegister_unitcell$3_9 VDDd out[5] Register_unitcell$3_9/q en default5 Register_unitcell$3_9/d
+ phi2 phi1 VSSd Register_unitcell$3
XRegister_unitcell$3_8 VDDd out[4] Register_unitcell$3_9/d en default4 Register_unitcell$3_8/d
+ phi2 phi1 VSSd Register_unitcell$3
.ends

.subckt scan_chain$1 VDDd ENd DATAd CLKd out[1] out[2] out[3] out[4] out[5] out[6]
+ out[7] out[8] out[9] out[10] out[20] out[19] out[18] out[17] out[16] out[15] out[14]
+ out[13] out[12] out[11] out[21] out[22] out[23] out[24] out[25] out[26] out[27]
+ out[28] out[29] out[30] out[40] out[39] out[38] out[37] out[36] out[35] out[34]
+ out[33] out[32] out[31] out[41] out[42] out[43] out[44] out[45] out[46] out[47]
+ out[48] out[49] out[50] VSSd
Xasc_hysteresis_buffer$9_0 VSSd CLKd VDDd SCHMITT$4_0/IN asc_hysteresis_buffer$9
Xasc_hysteresis_buffer$9_1 VSSd ENd VDDd SRegister_10$2_4/en asc_hysteresis_buffer$9
Xasc_hysteresis_buffer$9_2 VSSd DATAd VDDd SRegister_10$2_4/d asc_hysteresis_buffer$9
XSCHMITT$4_0 VDDd VSSd SCHMITT$4_0/IN SCHMITT$4_0/OUT SCHMITT$4
Xqw_NOLclk$2_0 SCHMITT$4_0/OUT VDDd VSSd qw_NOLclk$2_0/PHI_1 qw_NOLclk$2_0/PHI_2 qw_NOLclk$2
XSRegister_10$2_0 out[31] out[32] out[33] out[35] out[38] SRegister_10$2_3/q VSSd
+ VSSd VDDd VSSd VSSd VDDd VDDd VSSd VSSd VSSd out[39] out[36] out[34] out[40] SRegister_10$2_4/en
+ out[37] SRegister_10$2_2/d qw_NOLclk$2_0/PHI_2 VDDd VSSd qw_NOLclk$2_0/PHI_1 SRegister_10$2
XSRegister_10$2_2 out[41] out[42] out[43] out[45] out[48] SRegister_10$2_2/d VSSd
+ VSSd VSSd VSSd VDDd VSSd VSSd VDDd VDDd VSSd out[49] out[46] out[44] out[50] SRegister_10$2_4/en
+ out[47] SRegister_10$2_2/q qw_NOLclk$2_0/PHI_2 VDDd VSSd qw_NOLclk$2_0/PHI_1 SRegister_10$2
XSRegister_10$2_1 out[11] out[12] out[13] out[15] out[18] SRegister_10$2_4/q VSSd
+ VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd out[19] out[16] out[14] out[20] SRegister_10$2_4/en
+ out[17] SRegister_10$2_3/d qw_NOLclk$2_0/PHI_2 VDDd VSSd qw_NOLclk$2_0/PHI_1 SRegister_10$2
XSRegister_10$2_3 out[21] out[22] out[23] out[25] out[28] SRegister_10$2_3/d VSSd
+ VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd VSSd out[29] out[26] out[24] out[30] SRegister_10$2_4/en
+ out[27] SRegister_10$2_3/q qw_NOLclk$2_0/PHI_2 VDDd VSSd qw_NOLclk$2_0/PHI_1 SRegister_10$2
XSRegister_10$2_4 out[1] out[2] out[3] out[5] out[8] SRegister_10$2_4/d VSSd VSSd
+ VSSd VSSd VDDd VSSd VSSd VSSd VSSd VSSd out[9] out[6] out[4] out[10] SRegister_10$2_4/en
+ out[7] SRegister_10$2_4/q qw_NOLclk$2_0/PHI_2 VDDd VSSd qw_NOLclk$2_0/PHI_1 SRegister_10$2
.ends

.subckt pfet$457 a_254_0# a_348_560# w_n180_n88# a_414_0# a_n92_0# a_94_0# a_574_0#
+ a_508_560# a_188_560# a_28_560#
X0 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt pfet$455 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_348_n136# a_414_0#
+ a_n92_0# a_94_0# a_574_0# a_508_n136#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_n136# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_n136# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$484 a_254_0# a_350_460# a_414_0# a_n84_0# a_94_0# a_510_460# a_190_460#
+ a_574_0# a_30_460# VSUBS
X0 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_460# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_460# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt nfet$482 a_254_0# a_n84_0# a_94_0# a_190_460# a_30_460# VSUBS
X0 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$456 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
.ends

.subckt nfet$485 a_n84_0# a_94_0# a_30_460# VSUBS
X0 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt nfet$483 a_1054_0# a_734_0# a_254_0# a_350_460# a_830_460# a_894_0# a_990_460#
+ a_1214_0# a_414_0# a_n84_0# a_94_0# a_510_460# a_190_460# a_574_0# a_670_460# a_1150_460#
+ a_30_460# VSUBS
X0 a_734_0# a_670_460# a_574_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_574_0# a_510_460# a_414_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X3 a_1054_0# a_990_460# a_894_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X4 a_894_0# a_830_460# a_734_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X5 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X6 a_414_0# a_350_460# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X7 a_1214_0# a_1150_460# a_1054_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt Ncomparator$2 vss vdd out inn inp iref
Xpfet$457_1 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$457
Xpfet$457_2 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$457
Xpfet$455_0 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_570_1653# vdd m1_570_1653#
+ vdd m1_1242_549# pfet$455
Xpfet$457_3 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$457
Xpfet$455_1 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_1242_549# vdd m1_1242_549#
+ vdd m1_1242_549# pfet$455
Xpfet$455_3 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_1242_549# vdd m1_1242_549#
+ vdd m1_1242_549# pfet$455
Xpfet$455_2 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_570_1653# vdd m1_570_1653#
+ vdd m1_1242_549# pfet$455
Xnfet$484_0 vss iref m1_506_n191# vss m1_506_n191# iref iref vss iref vss nfet$484
Xnfet$484_1 vss iref iref vss iref iref iref vss iref vss nfet$484
Xnfet$484_2 m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191#
+ m1_506_n191# m1_506_n191# m1_506_n191# vss nfet$484
Xnfet$484_3 m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191#
+ m1_506_n191# m1_506_n191# m1_506_n191# vss nfet$484
Xnfet$482_0 m1_506_n191# m1_506_n191# m1_570_1653# inp inp vss nfet$482
Xnfet$484_5 vss iref m1_506_n191# vss m1_506_n191# iref iref vss iref vss nfet$484
Xnfet$484_4 vss iref iref vss iref iref iref vss iref vss nfet$484
Xnfet$482_1 m1_506_n191# m1_506_n191# m1_1242_549# inn inn vss nfet$482
Xnfet$482_3 m1_506_n191# m1_506_n191# m1_1242_549# inn inn vss nfet$482
Xnfet$482_2 m1_506_n191# m1_506_n191# m1_570_1653# inp inp vss nfet$482
Xpfet$456_0 vdd vdd vdd vdd vdd vdd pfet$456
Xpfet$456_1 vdd vdd vdd vdd vdd vdd pfet$456
Xpfet$456_2 vdd vdd vdd vdd vdd vdd pfet$456
Xpfet$456_3 vdd vdd vdd vdd vdd vdd pfet$456
Xnfet$485_1 vss vss vss vss nfet$485
Xnfet$485_0 vss vss vss vss nfet$485
Xnfet$483_0 out out vss iref iref vss iref vss out vss out iref iref vss iref iref
+ iref vss nfet$483
Xpfet$457_0 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$457
.ends

.subckt nfet$491 a_30_260# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_260# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$459 a_254_0# a_348_560# w_n180_n88# a_414_0# a_n92_0# a_94_0# a_574_0#
+ a_508_560# a_188_560# a_28_560#
X0 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$488 a_254_0# a_n84_0# a_94_0# a_190_460# a_30_460# VSUBS
X0 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt nfet$486 a_1054_0# a_734_0# a_510_n132# a_254_0# a_894_0# a_670_n132# a_1214_0#
+ a_830_n132# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132# a_574_0# a_990_n132#
+ a_350_n132# a_1150_n132# VSUBS
X0 a_734_0# a_670_n132# a_574_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X3 a_1054_0# a_990_n132# a_894_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X4 a_894_0# a_830_n132# a_734_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X5 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X6 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X7 a_1214_0# a_1150_n132# a_1054_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt pfet$460 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=1.625p ps=6.3u w=2.5u l=0.28u
.ends

.subckt pfet$458 a_1054_0# a_734_0# a_254_0# a_894_0# a_348_560# a_828_560# a_988_560#
+ w_n180_n88# a_1214_0# a_414_0# a_n92_0# a_94_0# a_574_0# a_508_560# a_188_560# a_668_560#
+ a_1148_560# a_28_560#
X0 a_1214_0# a_1148_560# a_1054_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_734_0# a_668_560# a_574_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X3 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X4 a_1054_0# a_988_560# a_894_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X5 a_894_0# a_828_560# a_734_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X6 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X7 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$487 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt Pcomparator$2 vss vdd out iref inn inp
Xpfet$459_4 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$459
Xpfet$459_6 vdd iref vdd iref vdd iref vdd iref iref iref pfet$459
Xpfet$459_5 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$459
Xnfet$488_0 vss vss m1_3615_n1223# m1_3615_n1223# m1_3615_n1223# vss nfet$488
Xpfet$459_7 vdd iref vdd iref vdd iref vdd iref iref iref pfet$459
Xnfet$488_1 vss vss m1_5539_n2811# m1_3615_n1223# m1_3615_n1223# vss nfet$488
Xpfet$459_8 vdd iref vdd iref vdd iref vdd iref iref iref pfet$459
Xnfet$488_2 vss vss m1_5539_n2811# m1_3615_n1223# m1_3615_n1223# vss nfet$488
Xnfet$486_0 out out m1_5539_n2811# vss vss m1_5539_n2811# vss m1_5539_n2811# out m1_5539_n2811#
+ vss out m1_5539_n2811# vss m1_5539_n2811# m1_5539_n2811# m1_5539_n2811# vss nfet$486
Xpfet$459_9 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$459
Xpfet$460_0 vdd vdd vdd vdd pfet$460
Xnfet$488_3 vss vss m1_3615_n1223# m1_3615_n1223# m1_3615_n1223# vss nfet$488
Xpfet$459_10 vdd iref vdd iref vdd iref vdd iref iref iref pfet$459
Xpfet$460_1 vdd vdd vdd vdd pfet$460
Xpfet$459_12 m1_2779_n1752# inn vdd m1_3615_n1223# m1_2779_n1752# m1_3615_n1223# m1_2779_n1752#
+ inn inn inn pfet$459
Xpfet$459_11 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$459
Xpfet$460_3 vdd vdd vdd vdd pfet$460
Xpfet$460_2 vdd vdd vdd vdd pfet$460
Xpfet$459_13 m1_2779_n1752# inp vdd m1_5539_n2811# m1_2779_n1752# m1_5539_n2811# m1_2779_n1752#
+ inp inp inp pfet$459
Xpfet$458_1 out out vdd vdd iref iref iref vdd vdd out vdd out vdd iref iref iref
+ iref iref pfet$458
Xpfet$458_0 out out vdd vdd iref iref iref vdd vdd out vdd out vdd iref iref iref
+ iref iref pfet$458
Xnfet$487_0 vss vss vss vss vss vss vss vss vss vss nfet$487
Xnfet$487_1 vss vss vss vss vss vss vss vss vss vss nfet$487
Xpfet$459_0 m1_2779_n1752# inp vdd m1_5539_n2811# m1_2779_n1752# m1_5539_n2811# m1_2779_n1752#
+ inp inp inp pfet$459
Xpfet$459_1 m1_2779_n1752# m1_2779_n1752# vdd m1_2779_n1752# m1_2779_n1752# m1_2779_n1752#
+ m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# pfet$459
Xpfet$459_2 m1_2779_n1752# inn vdd m1_3615_n1223# m1_2779_n1752# m1_3615_n1223# m1_2779_n1752#
+ inn inn inn pfet$459
Xpfet$459_3 m1_2779_n1752# m1_2779_n1752# vdd m1_2779_n1752# m1_2779_n1752# m1_2779_n1752#
+ m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# pfet$459
.ends

.subckt nfet$474 a_30_n132# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$450 a_28_460# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_460# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt nfet$479 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.5u
.ends

.subckt pfet$448 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# w_n180_n88# a_1262_n60# a_38_n60# a_n92_0# a_1058_n60# a_854_n60# a_342_0#
+ a_138_0# a_650_n60# a_1362_0#
X0 a_1362_0# a_1262_n60# a_1158_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X1 a_954_0# a_854_n60# a_750_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X2 a_1566_0# a_1466_n60# a_1362_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.5u
X3 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X4 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X5 a_1158_0# a_1058_n60# a_954_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X6 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.5u
X7 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
.ends

.subckt ppolyf_u_resistor$6 a_4000_0# a_n376_0# a_n132_0#
X0 a_n132_0# a_4000_0# a_n376_0# ppolyf_u r_width=1u r_length=20u
.ends

.subckt pfet$453 a_1054_0# a_734_0# a_828_n136# a_28_n136# a_254_0# a_894_0# a_188_n136#
+ a_988_n136# w_n180_n88# a_348_n136# a_1214_0# a_1148_n136# a_414_0# a_n92_0# a_94_0#
+ a_574_0# a_508_n136# a_668_n136#
X0 a_1214_0# a_1148_n136# a_1054_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_734_0# a_668_n136# a_574_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X3 a_574_0# a_508_n136# a_414_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X4 a_1054_0# a_988_n136# a_894_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X5 a_894_0# a_828_n136# a_734_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X6 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X7 a_414_0# a_348_n136# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt pfet$451 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$472 a_254_0# a_30_n132# a_n84_0# a_94_0# a_190_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$446 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_348_n136# a_414_0#
+ a_n92_0# a_94_0# a_574_0# a_508_n136#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_n136# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_n136# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$473 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt pfet$447 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
.ends

.subckt OTAforChargePump$3 vdd vss out iref inn inp
Xnfet$472_1 vss m1_116_n1334# vss m1_116_n1334# m1_116_n1334# vss nfet$472
Xnfet$472_2 vss m1_116_n1334# vss m1_116_n1334# m1_116_n1334# vss nfet$472
Xnfet$472_3 vss m1_116_n1334# vss out m1_116_n1334# vss nfet$472
Xpfet$446_1 inp m1_n400_n914# inp vdd inp m1_116_n1334# m1_n400_n914# m1_116_n1334#
+ m1_n400_n914# inp pfet$446
Xpfet$446_0 inn m1_n400_n914# inn vdd inn out m1_n400_n914# out m1_n400_n914# inn
+ pfet$446
Xpfet$446_2 iref vdd iref vdd iref iref vdd iref vdd iref pfet$446
Xpfet$446_3 iref vdd iref vdd iref m1_n400_n914# vdd m1_n400_n914# vdd iref pfet$446
Xpfet$446_4 iref vdd iref vdd iref m1_n400_n914# vdd m1_n400_n914# vdd iref pfet$446
Xpfet$446_5 iref vdd iref vdd iref iref vdd iref vdd iref pfet$446
Xpfet$446_6 iref vdd iref vdd iref iref vdd iref vdd iref pfet$446
Xpfet$446_7 iref vdd iref vdd iref m1_n400_n914# vdd m1_n400_n914# vdd iref pfet$446
Xpfet$446_8 inp m1_n400_n914# inp vdd inp m1_116_n1334# m1_n400_n914# m1_116_n1334#
+ m1_n400_n914# inp pfet$446
Xpfet$446_10 iref vdd iref vdd iref iref vdd iref vdd iref pfet$446
Xpfet$446_9 inn m1_n400_n914# inn vdd inn out m1_n400_n914# out m1_n400_n914# inn
+ pfet$446
Xnfet$473_1 vss vss vss vss vss vss vss vss vss vss nfet$473
Xnfet$473_0 vss vss vss vss vss vss vss vss vss vss nfet$473
Xpfet$446_11 iref vdd iref vdd iref m1_n400_n914# vdd m1_n400_n914# vdd iref pfet$446
Xpfet$447_0 m1_n400_n914# m1_n400_n914# m1_n400_n914# vdd m1_n400_n914# m1_n400_n914#
+ pfet$447
Xpfet$447_1 m1_n400_n914# m1_n400_n914# m1_n400_n914# vdd m1_n400_n914# m1_n400_n914#
+ pfet$447
Xpfet$447_2 vdd vdd vdd vdd vdd vdd pfet$447
Xpfet$447_3 vdd vdd vdd vdd vdd vdd pfet$447
Xpfet$447_4 vdd vdd vdd vdd vdd vdd pfet$447
Xpfet$447_5 vdd vdd vdd vdd vdd vdd pfet$447
Xnfet$472_0 vss m1_116_n1334# vss out m1_116_n1334# vss nfet$472
.ends

.subckt nfet$477 a_750_0# a_546_0# a_446_n132# a_n84_0# a_650_n132# a_38_n132# a_342_0#
+ a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_546_0# a_446_n132# a_342_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X2 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
X3 a_750_0# a_650_n132# a_546_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt nfet$475 a_750_0# a_546_0# a_446_n132# a_n84_0# a_650_n132# a_38_n132# a_342_0#
+ a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.5u
X1 a_546_0# a_446_n132# a_342_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.5u
X2 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.5u
X3 a_750_0# a_650_n132# a_546_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.5u
.ends

.subckt cap_mim$9 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=50u c_length=100u
.ends

.subckt nfet$480 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt pfet$449 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=0.8125p pd=3.8u as=0.325p ps=1.77u w=1.25u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.325p pd=1.77u as=0.8125p ps=3.8u w=1.25u l=0.5u
.ends

.subckt pfet$452 a_750_0# a_546_0# a_446_n60# a_242_n60# w_n180_n88# a_38_n60# a_n92_0#
+ a_342_0# a_138_0# a_650_n60#
X0 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X2 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.5u
.ends

.subckt nfet$478 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$476 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt PCP1248X$2 vdd s3 s2 s1 s0 vin iref200u out up down vss
Xnfet$474_4 m1_n539_12403# m1_16753_5552# vss vss nfet$474
Xpfet$450_8 m1_n539_12403# vdd OTAforChargePump$3_0/out m1_16753_5552# pfet$450
Xnfet$474_5 s0 OTAforChargePump$3_0/out m1_16753_5552# vss nfet$474
Xnfet$479_10 vss vss vss vss vss vss nfet$479
Xpfet$450_9 m1_n1311_12403# vdd OTAforChargePump$3_0/out m1_15009_5932# pfet$450
Xnfet$474_6 m1_n1311_12403# m1_15009_5932# vss vss nfet$474
Xnfet$479_11 vss vss vss vss vss vss nfet$479
Xpfet$448_30 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ pfet$448
Xnfet$474_7 s1 OTAforChargePump$3_0/out m1_15009_5932# vss nfet$474
Xppolyf_u_resistor$6_0 m1_3630_13790# vss m1_n502_13390# ppolyf_u_resistor$6
Xpfet$448_31 m1_n2925_n36# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187#
+ m1_1671_n1319# pfet$448
Xpfet$448_20 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ pfet$448
Xpfet$448_0 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$448
Xpfet$450_10 m1_n2083_12403# vdd OTAforChargePump$3_0/out m1_15881_3450# pfet$450
Xnfet$474_8 m1_n2083_12403# m1_15881_3450# vss vss nfet$474
Xppolyf_u_resistor$6_1 OTAforChargePump$3_0/inp vss m1_n502_13390# ppolyf_u_resistor$6
Xpfet$450_11 m1_n2855_12403# vdd OTAforChargePump$3_0/out m1_14137_3830# pfet$450
Xpfet$448_10 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$448
Xpfet$448_32 m1_n2925_n36# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187#
+ m1_1671_n1319# pfet$448
Xpfet$448_21 vdd vdd m1_1671_873# m1_1641_5849# m1_1641_5849# vdd m1_1671_873# m1_1641_5849#
+ vdd m1_1641_5849# m1_1641_5849# vdd m1_1641_5849# m1_1641_5849# vdd m1_1671_873#
+ m1_1641_5849# m1_1671_873# pfet$448
Xpfet$448_1 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$448
Xnfet$474_9 s2 OTAforChargePump$3_0/out m1_15881_3450# vss nfet$474
Xppolyf_u_resistor$6_2 m1_3630_14590# vss m1_n502_14190# ppolyf_u_resistor$6
Xpfet$448_11 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$448
Xpfet$448_22 vdd vdd m1_1671_n1319# m1_1137_12199# m1_1137_12199# vdd m1_1671_n1319#
+ m1_1137_12199# vdd m1_1137_12199# m1_1137_12199# vdd m1_1137_12199# m1_1137_12199#
+ vdd m1_1671_n1319# m1_1137_12199# m1_1671_n1319# pfet$448
Xpfet$448_33 vdd vdd m1_1671_n1319# m1_1137_12199# m1_1137_12199# vdd m1_1671_n1319#
+ m1_1137_12199# vdd m1_1137_12199# m1_1137_12199# vdd m1_1137_12199# m1_1137_12199#
+ vdd m1_1671_n1319# m1_1137_12199# m1_1671_n1319# pfet$448
Xpfet$448_2 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$448
Xpfet$453_0 m1_n2925_n36# m1_n2925_n36# up up out out up up vdd up out up m1_n2925_n36#
+ out m1_n2925_n36# out up up pfet$453
Xppolyf_u_resistor$6_3 m1_3630_13790# vss m1_n502_14190# ppolyf_u_resistor$6
Xnfet$479_0 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$479
Xpfet$448_12 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$448
Xpfet$448_23 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$448
Xpfet$448_34 vdd vdd m1_1671_n1319# m1_1137_12199# m1_1137_12199# vdd m1_1671_n1319#
+ m1_1137_12199# vdd m1_1137_12199# m1_1137_12199# vdd m1_1137_12199# m1_1137_12199#
+ vdd m1_1671_n1319# m1_1137_12199# m1_1671_n1319# pfet$448
Xpfet$448_3 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$448
Xppolyf_u_resistor$6_4 m1_3630_14590# vss m1_n502_14990# ppolyf_u_resistor$6
Xnfet$479_1 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$479
Xpfet$448_13 m1_n2925_n36# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187#
+ m1_1671_n1319# pfet$448
Xpfet$448_24 vdd vdd m1_n25_493# m1_n91_6229# m1_n91_6229# vdd m1_n25_493# m1_n91_6229#
+ vdd m1_n91_6229# m1_n91_6229# vdd m1_n91_6229# m1_n91_6229# vdd m1_n25_493# m1_n91_6229#
+ m1_n25_493# pfet$448
Xpfet$448_35 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ pfet$448
Xpfet$448_4 m1_n2925_n36# m1_n2925_n36# m1_n25_493# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n25_493# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36#
+ m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n25_493# m1_n1751_n2187# m1_n25_493#
+ pfet$448
Xppolyf_u_resistor$6_5 vdd vss m1_n502_14990# ppolyf_u_resistor$6
Xnfet$479_2 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$479
Xpfet$448_14 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$448
Xpfet$448_25 vdd vdd m1_1671_n1319# m1_1137_12199# m1_1137_12199# vdd m1_1671_n1319#
+ m1_1137_12199# vdd m1_1137_12199# m1_1137_12199# vdd m1_1137_12199# m1_1137_12199#
+ vdd m1_1671_n1319# m1_1137_12199# m1_1671_n1319# pfet$448
Xpfet$448_5 m1_n47_11059# m1_n47_11059# m1_6759_7857# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n47_11059# m1_6759_7857# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n47_11059# m1_n1751_n2187# m1_n1751_n2187# m1_n47_11059# m1_6759_7857# m1_n1751_n2187#
+ m1_6759_7857# pfet$448
Xpfet$451_0 vdd vdd m1_n2855_12403# s3 pfet$451
XOTAforChargePump$3_0 vdd vss OTAforChargePump$3_0/out iref200u vin OTAforChargePump$3_0/inp
+ OTAforChargePump$3
Xnfet$479_3 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$479
Xnfet$477_0 vss m1_9475_12045# OTAforChargePump$3_0/out vss OTAforChargePump$3_0/out
+ OTAforChargePump$3_0/out vss m1_9475_12045# OTAforChargePump$3_0/out vss nfet$477
Xpfet$448_6 vdd vdd m1_6759_7857# m1_n47_11059# m1_n47_11059# vdd m1_6759_7857# m1_n47_11059#
+ vdd m1_n47_11059# m1_n47_11059# vdd m1_n47_11059# m1_n47_11059# vdd m1_6759_7857#
+ m1_n47_11059# m1_6759_7857# pfet$448
Xpfet$448_15 m1_n2925_n36# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187#
+ m1_1671_n1319# pfet$448
Xpfet$448_26 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$448
Xpfet$451_1 vdd vdd m1_n2083_12403# s2 pfet$451
Xnfet$479_4 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$479
Xnfet$477_1 vss m1_n1751_n2187# OTAforChargePump$3_0/out vss OTAforChargePump$3_0/out
+ OTAforChargePump$3_0/out vss m1_n1751_n2187# OTAforChargePump$3_0/out vss nfet$477
Xpfet$448_7 vdd vdd m1_n25_493# m1_n91_6229# m1_n91_6229# vdd m1_n25_493# m1_n91_6229#
+ vdd m1_n91_6229# m1_n91_6229# vdd m1_n91_6229# m1_n91_6229# vdd m1_n25_493# m1_n91_6229#
+ m1_n25_493# pfet$448
Xpfet$448_16 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$448
Xpfet$448_27 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$448
Xpfet$451_2 vdd vdd m1_n539_12403# s0 pfet$451
Xnfet$479_5 m1_n47_11059# m1_n47_11059# m1_n47_11059# m1_n47_11059# m1_n47_11059#
+ vss nfet$479
Xnfet$477_2 vss m1_9475_12045# OTAforChargePump$3_0/out vss OTAforChargePump$3_0/out
+ OTAforChargePump$3_0/out vss m1_9475_12045# OTAforChargePump$3_0/out vss nfet$477
Xpfet$448_17 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$448
Xpfet$448_28 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ pfet$448
Xpfet$448_8 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$448
Xnfet$474_10 m1_n2855_12403# m1_14137_3830# vss vss nfet$474
Xpfet$451_3 vdd vdd m1_n1311_12403# s1 pfet$451
Xnfet$479_6 vss vss vss vss vss vss nfet$479
Xnfet$477_3 vss m1_n1751_n2187# OTAforChargePump$3_0/out vss OTAforChargePump$3_0/out
+ OTAforChargePump$3_0/out vss m1_n1751_n2187# OTAforChargePump$3_0/out vss nfet$477
Xpfet$448_18 m1_n2925_n36# m1_n2925_n36# m1_n25_493# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n25_493# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36#
+ m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n25_493# m1_n1751_n2187# m1_n25_493#
+ pfet$448
Xpfet$448_29 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$448
Xnfet$475_0 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$475
Xpfet$448_9 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$448
Xnfet$474_11 s3 OTAforChargePump$3_0/out m1_14137_3830# vss nfet$474
Xnfet$479_7 vss vss vss vss vss vss nfet$479
Xpfet$448_19 m1_n2925_n36# m1_n2925_n36# m1_1671_873# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_873# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36#
+ m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_873# m1_n1751_n2187# m1_1671_873#
+ pfet$448
Xnfet$475_1 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$475
Xnfet$479_8 vss vss vss vss vss vss nfet$479
Xcap_mim$9_0 m1_n1751_n2187# vdd cap_mim$9
Xnfet$475_2 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$475
Xnfet$480_0 down out m1_13543_n1758# down out m1_13543_n1758# down out down vss nfet$480
Xcap_mim$9_1 vss m1_9963_14448# cap_mim$9
Xnfet$479_9 vss vss vss vss vss vss nfet$479
Xnfet$475_3 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# vss nfet$475
Xcap_mim$9_2 vss OTAforChargePump$3_0/out cap_mim$9
Xnfet$475_4 m1_13543_n1758# m1_15039_784# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15039_784# m1_9963_14448# vss nfet$475
Xnfet$475_5 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# vss nfet$475
Xnfet$475_6 m1_13543_n1758# m1_16783_404# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_16783_404# m1_9963_14448# vss nfet$475
Xnfet$475_7 m1_13543_n1758# m1_15911_n1318# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15911_n1318# m1_9963_14448# vss nfet$475
Xpfet$449_0 vdd vdd vdd vdd vdd vdd pfet$449
Xnfet$475_8 m1_13543_n1758# m1_15911_n1318# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15911_n1318# m1_9963_14448# vss nfet$475
Xpfet$449_1 vdd vdd vdd m1_n1751_n2187# m1_n1751_n2187# m1_n1751_n2187# pfet$449
Xnfet$475_9 m1_13543_n1758# m1_15911_n1318# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15911_n1318# m1_9963_14448# vss nfet$475
Xpfet$449_2 vdd vdd vdd m1_9963_14448# m1_n1751_n2187# m1_n1751_n2187# pfet$449
Xnfet$475_30 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$475
Xpfet$449_3 vdd vdd vdd m1_n1751_n2187# m1_n1751_n2187# m1_n1751_n2187# pfet$449
Xnfet$475_20 vss m1_15911_n1318# m1_15881_3450# vss m1_15881_3450# m1_15881_3450#
+ vss m1_15911_n1318# m1_15881_3450# vss nfet$475
Xnfet$475_31 vss m1_14015_1164# OTAforChargePump$3_0/out vss OTAforChargePump$3_0/out
+ OTAforChargePump$3_0/out vss m1_14015_1164# OTAforChargePump$3_0/out vss nfet$475
Xpfet$449_4 vdd vdd vdd m1_9963_14448# m1_n1751_n2187# m1_n1751_n2187# pfet$449
Xnfet$475_21 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$475
Xnfet$475_32 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$475
Xnfet$475_10 m1_13543_n1758# m1_15911_n1318# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15911_n1318# m1_9963_14448# vss nfet$475
Xpfet$449_5 vdd vdd vdd vdd vdd vdd pfet$449
Xnfet$475_22 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$475
Xnfet$475_33 m1_n47_11059# m1_14015_1164# m1_9963_14448# m1_n47_11059# m1_9963_14448#
+ m1_9963_14448# m1_n47_11059# m1_14015_1164# m1_9963_14448# vss nfet$475
Xnfet$475_11 m1_13543_n1758# m1_15039_784# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15039_784# m1_9963_14448# vss nfet$475
Xpfet$452_0 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$452
Xnfet$478_0 s3 vss m1_n2855_12403# vss nfet$478
Xnfet$475_23 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$475
Xpfet$452_1 m1_n47_11059# m1_n47_11059# m1_n47_11059# m1_n47_11059# vdd m1_n47_11059#
+ m1_n47_11059# m1_n47_11059# m1_n47_11059# m1_n47_11059# pfet$452
Xnfet$475_34 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$475
Xnfet$475_12 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$475
Xnfet$478_1 s2 vss m1_n2083_12403# vss nfet$478
Xnfet$475_24 vss m1_15039_784# m1_15009_5932# vss m1_15009_5932# m1_15009_5932# vss
+ m1_15039_784# m1_15009_5932# vss nfet$475
Xnfet$475_35 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$475
Xpfet$452_2 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$452
Xnfet$475_13 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$475
Xnfet$478_2 s1 vss m1_n1311_12403# vss nfet$478
Xnfet$475_36 OTAforChargePump$3_0/inp m1_9475_12045# m1_9963_14448# OTAforChargePump$3_0/inp
+ m1_9963_14448# m1_9963_14448# OTAforChargePump$3_0/inp m1_9475_12045# m1_9963_14448#
+ vss nfet$475
Xnfet$475_25 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$475
Xpfet$452_3 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$452
Xpfet$452_10 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$452
Xnfet$475_14 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$475
Xpfet$450_0 m1_n539_12403# vdd m1_n47_11059# m1_1641_5849# pfet$450
Xnfet$478_3 s0 vss m1_n539_12403# vss nfet$478
Xnfet$476_0 vss vss vss vss vss vss nfet$476
Xpfet$452_11 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$452
Xnfet$475_26 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$475
Xnfet$475_15 vss vss vss vss vss vss vss vss vss vss nfet$475
Xpfet$452_4 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$452
Xpfet$450_1 s0 vdd m1_1641_5849# vdd pfet$450
Xnfet$476_1 vss vss vss vss vss vss nfet$476
Xnfet$475_27 vss m1_15911_n1318# m1_15881_3450# vss m1_15881_3450# m1_15881_3450#
+ vss m1_15911_n1318# m1_15881_3450# vss nfet$475
Xnfet$475_16 vss vss vss vss vss vss vss vss vss vss nfet$475
Xpfet$452_5 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$452
Xpfet$450_2 s3 vdd m1_n1771_4009# vdd pfet$450
Xnfet$476_2 vss m1_9963_14448# vss m1_9963_14448# m1_9963_14448# vss nfet$476
Xnfet$475_28 vss m1_15911_n1318# m1_15881_3450# vss m1_15881_3450# m1_15881_3450#
+ vss m1_15911_n1318# m1_15881_3450# vss nfet$475
Xnfet$475_17 vss m1_16783_404# m1_16753_5552# vss m1_16753_5552# m1_16753_5552# vss
+ m1_16783_404# m1_16753_5552# vss nfet$475
Xpfet$452_6 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$452
Xpfet$450_3 m1_n1311_12403# vdd m1_n47_11059# m1_n91_6229# pfet$450
Xnfet$475_29 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$475
Xnfet$475_18 vss m1_15039_784# m1_15009_5932# vss m1_15009_5932# m1_15009_5932# vss
+ m1_15039_784# m1_15009_5932# vss nfet$475
Xnfet$474_0 s0 m1_n47_11059# m1_1641_5849# vss nfet$474
Xpfet$452_7 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$452
Xpfet$450_4 m1_n2083_12403# vdd m1_n47_11059# m1_1137_12199# pfet$450
Xnfet$475_19 vss m1_15911_n1318# m1_15881_3450# vss m1_15881_3450# m1_15881_3450#
+ vss m1_15911_n1318# m1_15881_3450# vss nfet$475
Xpfet$452_8 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$452
Xnfet$474_1 s1 m1_n47_11059# m1_n91_6229# vss nfet$474
Xpfet$450_5 m1_n2855_12403# vdd m1_n47_11059# m1_n1771_4009# pfet$450
Xnfet$474_2 s3 m1_n47_11059# m1_n1771_4009# vss nfet$474
Xpfet$452_9 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$452
Xpfet$450_6 s1 vdd m1_n91_6229# vdd pfet$450
Xnfet$474_3 s2 m1_n47_11059# m1_1137_12199# vss nfet$474
Xpfet$450_7 s2 vdd m1_1137_12199# vdd pfet$450
.ends

.subckt pfet$463 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt ppolyf_u_resistor$7 a_n376_0# a_4200_0# a_n132_0#
X0 a_n132_0# a_4200_0# a_n376_0# ppolyf_u r_width=1u r_length=21u
.ends

.subckt cap_mim$10 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=60u c_length=100u
.ends

.subckt pfet$462 a_28_460# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_460# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt nfet$489 a_n84_0# a_94_0# a_30_460# VSUBS
X0 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$461 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=2.6p pd=9.3u as=2.6p ps=9.3u w=4u l=0.28u
.ends

.subckt nfet$490 a_30_n132# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt SCHMITT$5 VDD VSS IN OUT
Xpfet$462_0 OUT VDD m1_596_1544# VSS pfet$462
Xnfet$489_0 m1_592_402# OUT IN VSS nfet$489
Xnfet$489_1 VSS m1_592_402# IN VSS nfet$489
Xpfet$461_0 IN VDD m1_596_1544# OUT pfet$461
Xpfet$461_1 IN VDD VDD m1_596_1544# pfet$461
Xnfet$490_0 OUT m1_592_402# VDD VSS nfet$490
.ends

.subckt pfet$454 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt nfet$481 a_n84_0# a_94_0# a_30_160# VSUBS
X0 a_94_0# a_30_160# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.28u
.ends

.subckt SRLATCH$1 vdd vss q qb s r
Xpfet$454_0 r vdd m1_818_875# qb pfet$454
Xpfet$454_1 q vdd vdd m1_818_875# pfet$454
Xpfet$454_2 s vdd m1_50_875# vdd pfet$454
Xpfet$454_3 qb vdd q m1_50_875# pfet$454
Xnfet$481_0 vss qb r vss nfet$481
Xnfet$481_1 vss qb q vss nfet$481
Xnfet$481_2 q vss s vss nfet$481
Xnfet$481_3 q vss qb vss nfet$481
.ends

.subckt VCOfinal$1 s3 s0 s1 s2 iref200 fout foutb irefp irefn vin a_11641_n18839#
+ vdd vss
XNcomparator$2_0 vss vdd SRLATCH$1_0/s Ncomparator$2_0/inn PCP1248X$2_0/out irefn
+ Ncomparator$2
Xnfet$491_0 SRLATCH$1_0/q vss PCP1248X$2_0/up vss nfet$491
Xnfet$491_1 SCHMITT$5_0/OUT vss foutb vss nfet$491
Xnfet$491_2 SCHMITT$5_1/OUT vss fout vss nfet$491
XPcomparator$2_0 vss vdd SRLATCH$1_0/r irefp PCP1248X$2_0/out Pcomparator$2_0/inp
+ Pcomparator$2
XPCP1248X$2_0 vdd s3 s2 s1 s0 vin iref200 PCP1248X$2_0/out PCP1248X$2_0/up SRLATCH$1_0/qb
+ vss PCP1248X$2
Xpfet$463_0 SRLATCH$1_0/q vdd vdd PCP1248X$2_0/up pfet$463
Xpfet$463_1 SCHMITT$5_0/OUT vdd vdd foutb pfet$463
Xpfet$463_2 SCHMITT$5_1/OUT vdd vdd fout pfet$463
Xppolyf_u_resistor$7_0 vss vss Pcomparator$2_0/inp ppolyf_u_resistor$7
Xppolyf_u_resistor$7_1 vss m1_13996_n13334# Ncomparator$2_0/inn ppolyf_u_resistor$7
Xppolyf_u_resistor$7_2 vss m1_13996_n13334# Pcomparator$2_0/inp ppolyf_u_resistor$7
Xppolyf_u_resistor$7_3 vss vdd Ncomparator$2_0/inn ppolyf_u_resistor$7
Xcap_mim$10_0 vss PCP1248X$2_0/out cap_mim$10
XSCHMITT$5_0 vdd vss SRLATCH$1_0/qb SCHMITT$5_0/OUT SCHMITT$5
XSCHMITT$5_1 vdd vss SRLATCH$1_0/q SCHMITT$5_1/OUT SCHMITT$5
XSRLATCH$1_0 vdd vss SRLATCH$1_0/q SRLATCH$1_0/qb SRLATCH$1_0/s SRLATCH$1_0/r SRLATCH$1
.ends

.subckt nfet$433 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$407 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$432 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$408 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt xp_3_1_MUX$5 S0 S1 VDD VSS OUT_1 C_1 B_1 A_1
Xnfet$433_0 S1 VSS m1_n432_n1290# VSS nfet$433
Xnfet$433_1 S0 VSS m1_n432_458# VSS nfet$433
Xpfet$407_0 VDD A_1 m1_239_n318# m1_n432_458# pfet$407
Xpfet$407_2 VDD B_1 m1_239_n318# S0 pfet$407
Xpfet$407_1 VDD C_1 OUT_1 S1 pfet$407
Xpfet$407_3 VDD m1_239_n318# OUT_1 m1_n432_n1290# pfet$407
Xnfet$432_0 m1_n432_n1290# C_1 OUT_1 VSS nfet$432
Xnfet$432_1 m1_n432_458# B_1 m1_239_n318# VSS nfet$432
Xnfet$432_2 S1 m1_239_n318# OUT_1 VSS nfet$432
Xnfet$432_3 S0 A_1 m1_239_n318# VSS nfet$432
Xpfet$408_0 VDD VDD m1_n432_n1290# S1 pfet$408
Xpfet$408_1 VDD VDD m1_n432_458# S0 pfet$408
.ends

.subckt pfet$356 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$349 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$371 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$378 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$351 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$389 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$354 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$375 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$352 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$396 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$372 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$392 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$377 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$397 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$390 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$375 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$403 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$348 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$383 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$368 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$370 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$350 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$373 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$376 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$380 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$369 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$373 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$401 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$374 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$399 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$381 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$366 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$359 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$374 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$371 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$364 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$357 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$395 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$362 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$388 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$355 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$393 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$378 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$353 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$360 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$386 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$379 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$391 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$376 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$404 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$384 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$369 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$377 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$402 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$367 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$382 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$372 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$400 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$398 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$380 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$365 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$358 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$370 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$363 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$394 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$379 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$361 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$387 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$405 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$385 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_dual_psd_def_20250809$5 vdd vss pd1 pd2 pd3 pd4 pd5 pd6 pd7 pd8 pd9 fout
+ sd1 sd2 sd3 sd4 sd5 sd6 sd7 sd8 sd9 fin define
Xpfet$356_6 vdd vdd m1_n290_24224# m1_n910_23922# pfet$356
Xpfet$349_5 vdd m1_7198_15778# m1_6377_16202# m1_6116_17343# pfet$349
Xnfet$371_6 m1_2384_21590# m1_2384_21590# m1_3871_22513# m1_3871_22513# m1_2843_21586#
+ vss nfet$371
Xnfet$378_10 m1_32675_25947# vss m1_35071_24542# vss nfet$378
Xpfet$351_19 vdd m1_n3822_20130# m1_n3822_20130# m1_27441_19850# m1_27003_19550# m1_27003_19550#
+ pfet$351
Xnfet$389_20 m1_22493_16080# m1_22493_16080# m1_22034_17714# m1_22034_17714# m1_22591_16398#
+ vss nfet$389
Xpfet$354_3 vdd vdd m1_5901_19550# m1_649_17714# pfet$354
Xnfet$375_11 m1_9331_15478# vss m1_15171_20152# vss nfet$375
Xpfet$352_0 vdd vdd m1_n1133_21590# m1_n1263_21786# pfet$352
Xnfet$389_7 m1_5761_16080# m1_5761_16080# m1_5302_17714# m1_5302_17714# m1_5859_16398#
+ vss nfet$389
Xnfet$396_8 m1_9624_19404# m1_9624_19404# vss vss m1_n3724_21430# vss nfet$396
Xpfet$349_108 vdd vdd m1_15454_18030# m1_15564_15778# pfet$349
Xnfet$372_12 m1_16452_19550# m1_16452_19550# vss vss m1_16890_20470# vss nfet$372
Xnfet$392_2 m1_n6274_17836# m1_n5351_15778# m1_n6172_16202# vss nfet$392
Xnfet$378_0 m1_n10452_25858# vss m1_n1271_25858# vss nfet$378
Xpfet$349_19 vdd m1_3015_15778# m1_2194_16202# m1_1933_17343# pfet$349
Xpfet$377_2 vdd m1_n5764_21786# m1_n5764_21786# m1_n5019_22344# m1_n5227_21418# m1_n5227_21418#
+ pfet$377
Xnfet$371_7 m1_5771_21786# m1_5771_21786# m1_7388_22513# m1_7388_22513# m1_6992_21586#
+ vss nfet$371
Xnfet$378_11 m1_32554_23922# vss m1_33174_24224# vss nfet$378
Xpfet$356_7 vdd vdd m1_32330_25662# m1_32193_25858# pfet$356
Xpfet$349_6 vdd vdd m1_7198_15778# m1_7555_16080# pfet$349
Xnfet$389_21 m1_14127_16080# m1_14127_16080# vss vss m1_15690_17358# vss nfet$389
Xnfet$389_10 m1_1578_16080# m1_1578_16080# m1_1119_17714# m1_1119_17714# m1_1676_16398#
+ vss nfet$389
Xpfet$354_4 vdd vdd m1_12935_19550# m1_9015_17714# pfet$354
Xnfet$375_12 m1_13514_15478# vss m1_18688_20152# vss nfet$375
Xpfet$352_1 vdd vdd m1_11671_21786# m1_11039_21786# pfet$352
Xnfet$389_8 m1_3015_15778# m1_3015_15778# m1_2905_18030# m1_2905_18030# m1_3141_17358#
+ vss nfet$389
Xnfet$396_9 m1_n6380_21786# m1_n6380_21786# m1_n6839_21786# m1_n6839_21786# m1_n6282_21430#
+ vss nfet$396
Xpfet$349_109 vdd vdd m1_10299_17343# m1_13198_17714# pfet$349
Xnfet$372_13 m1_19969_19550# m1_19969_19550# vss vss m1_20407_20470# vss nfet$372
Xnfet$397_10 vss vss m1_n4978_24224# vss nfet$397
Xnfet$392_3 m1_n6433_17343# m1_n6172_16202# m1_n6657_17518# vss nfet$392
Xnfet$378_1 m1_n789_25858# vss m1_n647_25662# vss nfet$378
Xnfet$371_8 m1_23486_21590# m1_23486_21590# m1_24973_22513# m1_24973_22513# m1_23945_21586#
+ vss nfet$371
Xnfet$378_12 m1_32675_25947# vss m1_28624_21786# vss nfet$378
Xpfet$356_8 vdd vdd m1_33174_24224# m1_32554_23922# pfet$356
Xnfet$390_0 m1_4620_20152# m1_4620_20152# m1_2590_19404# m1_2590_19404# m1_3454_20470#
+ vss nfet$390
Xpfet$349_7 vdd vdd m1_6275_17836# m1_6116_17343# pfet$349
Xpfet$375_0 vdd vdd m1_n7186_25858# m1_n10452_25858# pfet$375
Xpfet$354_5 vdd vdd m1_8137_20152# m1_965_15478# pfet$354
Xnfet$403_0 m1_n927_19404# m1_n927_19404# vss vss m1_n6282_20470# vss nfet$403
Xnfet$389_22 m1_15564_15778# m1_15564_15778# m1_15454_18030# m1_15454_18030# m1_15690_17358#
+ vss nfet$389
Xnfet$389_11 m1_6377_16202# m1_6377_16202# vss vss m1_5859_16398# vss nfet$389
Xnfet$375_13 m1_13198_17714# vss m1_16452_19550# vss nfet$375
Xpfet$352_2 vdd vdd m1_12935_21590# m1_12805_21786# pfet$352
Xnfet$389_9 m1_2194_16202# m1_2194_16202# vss vss m1_1676_16398# vss nfet$389
Xpfet$348_110 vdd m1_11903_24542# vdd m1_12875_24346# pfet$348
Xnfet$372_14 m1_17381_17714# m1_17381_17714# vss vss m1_21039_20470# vss nfet$372
Xnfet$397_11 m1_n10452_25858# vss m1_n4847_25662# vss nfet$397
Xnfet$392_4 m1_27031_17343# m1_27292_16202# m1_26807_17518# vss nfet$392
Xnfet$378_2 m1_n1271_25858# vss m1_n1134_25662# vss nfet$378
Xnfet$371_9 m1_23356_21786# m1_23356_21786# m1_24973_22513# m1_24973_22513# m1_24577_21586#
+ vss nfet$371
Xnfet$378_13 m1_32675_25947# vss m1_32817_25662# vss nfet$378
Xpfet$356_9 vdd vdd m1_28624_21786# m1_32675_25947# pfet$356
Xnfet$383_0 m1_21456_22513# m1_21456_22513# m1_30256_19792# m1_30256_19792# m1_30492_20470#
+ vss nfet$383
Xnfet$390_1 m1_1103_20152# m1_1103_20152# m1_n927_19404# m1_n927_19404# m1_n63_20470#
+ vss nfet$390
Xpfet$349_8 vdd vdd m1_9331_15478# sd5 pfet$349
Xpfet$368_0 vdd vdd m1_n7513_20152# m1_35837_22102# pfet$368
Xpfet$375_1 vdd m1_n7186_25858# vdd m1_n6111_25858# pfet$375
Xnfet$403_1 m1_n2543_20130# m1_n2543_20130# m1_n5227_20152# m1_n5227_20152# m1_n2445_20470#
+ vss nfet$403
Xnfet$389_23 m1_18926_16202# m1_18926_16202# vss vss m1_18408_16398# vss nfet$389
Xpfet$354_6 vdd vdd m1_9418_19550# m1_4832_17714# pfet$354
Xnfet$389_12 m1_n1168_15778# m1_n1168_15778# m1_n1278_18030# m1_n1278_18030# m1_n1042_17358#
+ vss nfet$389
Xnfet$370_80 m1_28147_25662# m1_28991_24224# m1_30095_25658# vss nfet$370
Xpfet$352_10 vdd vdd m1_23486_21590# m1_23356_21786# pfet$352
Xnfet$375_14 m1_21564_17714# vss m1_23486_19550# vss nfet$375
Xpfet$352_3 vdd vdd m1_9418_21590# m1_9288_21786# pfet$352
Xpfet$348_100 vdd vdd m1_29607_24346# m1_n7513_20152# pfet$348
Xpfet$350_0 vdd vdd vdd m1_n674_22102# m1_n1133_21590# m1_n1133_21590# pfet$350
Xnfet$372_15 m1_21564_17714# m1_21564_17714# vss vss m1_24556_20470# vss nfet$372
Xnfet$397_12 m1_n10452_25858# vss m1_n5571_25662# vss nfet$397
Xnfet$392_5 m1_27031_17343# m1_29087_15778# m1_28470_16080# vss nfet$392
Xnfet$378_3 m1_n7513_20152# vss m1_326_24346# vss nfet$378
Xnfet$373_80 m1_18824_17836# m1_19747_15778# m1_18926_16202# vss nfet$373
Xnfet$383_1 m1_14422_22513# m1_14422_22513# m1_31535_19792# m1_31535_19792# m1_31771_20470#
+ vss nfet$383
Xnfet$390_2 m1_n3218_15478# m1_n3218_15478# m1_2590_19404# m1_2590_19404# m1_2822_20470#
+ vss nfet$390
Xpfet$349_9 vdd vdd m1_8172_15778# m1_5302_17714# pfet$349
Xnfet$376_0 sd9 vss m1_n7401_15478# vss nfet$376
Xnfet$389_24 m1_18310_16080# m1_18310_16080# m1_17851_17714# m1_17851_17714# m1_18408_16398#
+ vss nfet$389
Xpfet$354_7 vdd vdd m1_11654_20152# m1_5148_15478# pfet$354
Xnfet$389_13 m1_n2605_16080# m1_n2605_16080# vss vss m1_n1042_17358# vss nfet$389
Xnfet$370_81 m1_n7513_20152# vss m1_25424_24346# vss nfet$370
Xnfet$370_70 m1_21590_21786# vss m1_28010_25858# vss nfet$370
Xpfet$352_11 vdd vdd m1_18705_21786# m1_18073_21786# pfet$352
Xpfet$380_0 vdd vdd m1_n8145_21908# m1_n6839_20152# pfet$380
Xnfet$375_15 m1_17697_15478# vss m1_22205_20152# vss nfet$375
Xpfet$352_4 vdd vdd m1_8154_21786# m1_7522_21786# pfet$352
Xpfet$350_1 vdd m1_7388_22513# m1_7388_22513# m1_6988_22402# m1_7522_21786# m1_7522_21786#
+ pfet$350
Xpfet$348_101 vdd vdd m1_28010_25858# m1_21590_21786# pfet$348
Xnfet$372_16 m1_23486_19550# m1_23486_19550# vss vss m1_23924_20470# vss nfet$372
Xnfet$397_13 fin vss m1_n4623_25487# vss nfet$397
Xnfet$392_6 m1_27190_17836# m1_28113_15778# m1_27292_16202# vss nfet$392
Xnfet$378_4 m1_n789_25858# vss m1_1607_24542# vss nfet$378
Xnfet$373_81 m1_13198_17714# vss m1_10299_17343# vss nfet$373
Xnfet$373_70 m1_n7513_20152# vss m1_18310_16080# vss nfet$373
Xnfet$376_1 sd2 vss m1_21880_15478# vss nfet$376
Xnfet$383_2 m1_17939_22513# m1_17939_22513# vss vss m1_31771_20470# vss nfet$383
Xnfet$390_3 m1_8137_20152# m1_8137_20152# m1_6107_19404# m1_6107_19404# m1_6971_20470#
+ vss nfet$390
Xnfet$369_0 m1_4509_24346# m1_4509_24346# vss vss m1_3991_24542# vss nfet$369
Xnfet$389_25 m1_14743_16202# m1_14743_16202# vss vss m1_14225_16398# vss nfet$389
Xnfet$389_14 m1_n2605_16080# m1_n2605_16080# m1_n3064_17714# m1_n3064_17714# m1_n2507_16398#
+ vss nfet$389
Xpfet$354_8 vdd vdd m1_n1133_19550# m1_n7383_17599# pfet$354
Xnfet$370_82 m1_11415_25662# m1_12259_24224# m1_13363_25658# vss nfet$370
Xnfet$370_71 m1_28147_25662# m1_28371_23922# m1_28635_24542# vss nfet$370
Xnfet$370_60 pd6 vss m1_16322_21786# vss nfet$370
Xpfet$352_12 vdd vdd m1_16452_21590# m1_16322_21786# pfet$352
Xpfet$373_0 vdd vdd m1_n4485_20152# m1_n3822_20130# pfet$373
Xnfet$375_16 m1_17381_17714# vss m1_19969_19550# vss nfet$375
Xnfet$401_0 m1_n8283_20611# vss m1_n8283_19850# vss nfet$401
Xpfet$352_5 vdd vdd m1_1120_21786# m1_488_21786# pfet$352
Xpfet$350_2 vdd m1_7388_22513# m1_7388_22513# m1_6360_22102# m1_8154_21786# m1_8154_21786#
+ pfet$350
Xpfet$348_102 vdd m1_28371_23922# m1_28635_24542# m1_28010_25858# pfet$348
Xpfet$374_10 vdd vdd m1_n10933_25858# fin pfet$374
Xnfet$372_17 m1_12935_19550# m1_12935_19550# vss vss m1_13373_20470# vss nfet$372
Xnfet$399_0 m1_n10933_25858# m1_n8848_25658# m1_n8055_24542# vss nfet$399
Xnfet$392_7 m1_27190_17836# m1_28470_16080# m1_28003_18030# vss nfet$392
Xnfet$378_5 m1_n789_25858# vss m1_488_21786# vss nfet$378
Xnfet$373_82 m1_10299_17343# vss m1_10458_17836# vss nfet$373
Xnfet$373_71 m1_14641_17836# m1_15921_16080# m1_15454_18030# vss nfet$373
Xnfet$373_60 m1_18665_17343# vss m1_18824_17836# vss nfet$373
Xnfet$376_2 sd1 vss m1_26063_15478# vss nfet$376
Xnfet$383_3 m1_24973_22513# m1_24973_22513# vss vss m1_30492_20470# vss nfet$383
Xnfet$390_4 m1_965_15478# m1_965_15478# m1_6107_19404# m1_6107_19404# m1_6339_20470#
+ vss nfet$390
Xnfet$369_1 m1_3893_24224# m1_3893_24224# m1_3537_24542# m1_3537_24542# m1_3991_24542#
+ vss nfet$369
Xnfet$389_26 m1_14127_16080# m1_14127_16080# m1_13668_17714# m1_13668_17714# m1_14225_16398#
+ vss nfet$389
Xpfet$354_9 vdd vdd m1_27003_19550# m1_25747_17714# pfet$354
Xnfet$389_15 m1_n1989_16202# m1_n1989_16202# vss vss m1_n2507_16398# vss nfet$389
Xnfet$381_0 m1_n290_24224# m1_n290_24224# m1_n646_24542# m1_n646_24542# m1_n192_24542#
+ vss nfet$381
Xnfet$370_72 m1_23827_25858# m1_25912_25658# m1_26705_24542# vss nfet$370
Xnfet$370_61 m1_23964_25662# m1_24808_24224# m1_25912_25658# vss nfet$370
Xnfet$370_50 m1_n7513_20152# vss m1_21241_24346# vss nfet$370
Xpfet$352_13 vdd vdd m1_15188_21786# m1_14556_21786# pfet$352
Xpfet$366_0 vdd vdd m1_n7247_17714# m1_n6788_16080# pfet$366
Xpfet$373_1 vdd m1_n4485_21904# vdd m1_9624_19404# pfet$373
Xnfet$375_17 m1_21880_15478# vss m1_25722_20152# vss nfet$375
Xnfet$401_1 m1_n7513_20152# m1_n8283_19850# vss vss nfet$401
Xpfet$352_6 vdd vdd m1_5901_21590# m1_5771_21786# pfet$352
Xpfet$348_103 vdd vdd m1_28635_24542# m1_28991_24224# pfet$348
Xpfet$350_3 vdd m1_9645_21447# m1_9645_21447# m1_10505_22402# m1_11039_21786# m1_11039_21786#
+ pfet$350
Xnfet$399_1 m1_n10796_25662# m1_n10572_23922# m1_n10308_24542# vss nfet$399
Xpfet$374_11 vdd vdd m1_n9336_24346# vss pfet$374
Xnfet$378_6 m1_n910_23922# vss m1_n290_24224# vss nfet$378
Xnfet$373_72 m1_17851_17714# vss m1_18441_17518# vss nfet$373
Xnfet$373_61 m1_20104_16080# vss m1_19747_15778# vss nfet$373
Xnfet$373_50 m1_25747_17714# vss m1_22848_17343# vss nfet$373
Xnfet$383_4 m1_32818_20470# m1_32818_20470# vss vss m1_34329_20470# vss nfet$383
Xnfet$369_2 m1_4997_25658# m1_4997_25658# vss vss m1_5456_25502# vss nfet$369
Xnfet$390_5 m1_5148_15478# m1_5148_15478# m1_9624_19404# m1_9624_19404# m1_9856_20470#
+ vss nfet$390
Xnfet$381_1 m1_814_25658# m1_814_25658# vss vss m1_1273_25502# vss nfet$381
Xnfet$370_73 m1_24309_25858# vss m1_21590_21786# vss nfet$370
Xnfet$370_62 m1_24188_23922# vss m1_24808_24224# vss nfet$370
Xnfet$370_51 m1_19644_25858# m1_21729_25658# m1_22522_24542# vss nfet$370
Xnfet$370_40 m1_15598_25662# m1_16442_24224# m1_17546_25658# vss nfet$370
Xnfet$389_27 m1_18310_16080# m1_18310_16080# vss vss m1_19873_17358# vss nfet$389
Xnfet$389_16 m1_19747_15778# m1_19747_15778# m1_19637_18030# m1_19637_18030# m1_19873_17358#
+ vss nfet$389
Xpfet$359_0 vdd m1_31535_19792# vdd m1_17939_22513# pfet$359
Xpfet$366_1 vdd m1_n7247_17714# vdd m1_n6172_16202# pfet$366
Xnfet$374_0 m1_n1263_21786# vss m1_n1133_21590# vss nfet$374
Xpfet$373_2 vdd m1_n5227_21418# vdd m1_2590_19404# pfet$373
Xpfet$352_14 vdd vdd m1_19969_21590# m1_19839_21786# pfet$352
Xnfet$401_2 m1_n8145_21908# vss m1_n8283_20611# vss nfet$401
Xpfet$352_7 vdd vdd m1_4637_21786# m1_4005_21786# pfet$352
Xpfet$348_104 vdd m1_25912_25658# m1_26705_24542# m1_23964_25662# pfet$348
Xpfet$350_4 vdd vdd vdd m1_9877_22102# m1_9418_21590# m1_9418_21590# pfet$350
Xnfet$399_2 m1_n10933_25858# m1_n10309_25662# m1_n10572_23922# vss nfet$399
Xpfet$374_12 vdd vdd m1_n7082_23622# m1_n8625_26174# pfet$374
Xpfet$348_90 vdd vdd m1_24309_25858# m1_25424_24346# pfet$348
Xnfet$378_7 m1_25107_21786# vss m1_32193_25858# vss nfet$378
Xnfet$373_73 m1_13668_17714# vss m1_16538_15778# vss nfet$373
Xnfet$373_62 m1_18665_17343# m1_20721_15778# m1_20104_16080# vss nfet$373
Xnfet$373_51 m1_n7513_20152# vss m1_22493_16080# vss nfet$373
Xnfet$373_40 m1_n2250_17343# m1_n194_15778# m1_n811_16080# vss nfet$373
Xnfet$383_5 m1_32818_21586# m1_32818_21586# m1_34093_19792# m1_34093_19792# m1_34329_20470#
+ vss nfet$383
Xnfet$369_3 m1_4509_24346# m1_4509_24346# m1_3394_25858# m1_3394_25858# m1_5456_25502#
+ vss nfet$369
Xnfet$390_6 m1_11654_20152# m1_11654_20152# m1_9624_19404# m1_9624_19404# m1_10488_20470#
+ vss nfet$390
Xnfet$370_52 m1_20126_25858# vss m1_22522_24542# vss nfet$370
Xnfet$370_41 pd5 vss m1_12805_21786# vss nfet$370
Xnfet$370_30 m1_n7513_20152# vss m1_17058_24346# vss nfet$370
Xnfet$389_17 m1_22493_16080# m1_22493_16080# vss vss m1_24056_17358# vss nfet$389
Xnfet$381_2 m1_326_24346# m1_326_24346# m1_n789_25858# m1_n789_25858# m1_1273_25502#
+ vss nfet$381
Xpfet$366_2 vdd vdd m1_n5461_18030# m1_n5351_15778# pfet$366
Xpfet$373_3 vdd vdd m1_n5227_21418# m1_6107_19404# pfet$373
Xnfet$374_1 m1_11039_21786# vss m1_11671_21786# vss nfet$374
Xnfet$370_74 pd8 vss m1_23356_21786# vss nfet$370
Xpfet$352_15 vdd vdd m1_27003_21590# m1_26873_21786# pfet$352
Xnfet$370_63 m1_14556_21786# vss m1_19644_25858# vss nfet$370
Xpfet$359_1 vdd vdd m1_30256_19792# m1_21456_22513# pfet$359
Xnfet$401_3 m1_n8283_19850# m1_n8283_20611# vss vss nfet$401
Xpfet$352_8 vdd vdd m1_2384_21590# m1_2254_21786# pfet$352
Xpfet$371_0 vdd vdd m1_n7320_25516# m1_n7186_25858# pfet$371
Xpfet$348_105 vdd vdd m1_30888_24542# m1_28492_25858# pfet$348
Xpfet$350_5 vdd m1_9645_21447# m1_9645_21447# m1_9877_22102# m1_11671_21786# m1_11671_21786#
+ pfet$350
Xpfet$374_13 vdd vdd m1_n8055_24542# m1_n8625_26174# pfet$374
Xpfet$348_91 vdd vdd m1_23356_21786# pd8 pfet$348
Xpfet$348_80 vdd vdd m1_17058_24346# m1_n7513_20152# pfet$348
Xnfet$399_3 m1_n10796_25662# m1_n9952_24224# m1_n8848_25658# vss nfet$399
Xnfet$378_8 m1_32193_25858# vss m1_32330_25662# vss nfet$378
Xnfet$397_0 m1_n8625_26174# vss m1_n8055_24542# vss nfet$397
Xnfet$373_74 m1_14482_17343# vss m1_14641_17836# vss nfet$373
Xnfet$373_63 m1_13668_17714# vss m1_14258_17518# vss nfet$373
Xnfet$373_52 m1_23007_17836# m1_24287_16080# m1_23820_18030# vss nfet$373
Xnfet$373_30 sd6 vss m1_5148_15478# vss nfet$373
Xnfet$373_41 m1_n2091_17836# m1_n1168_15778# m1_n1989_16202# vss nfet$373
Xnfet$383_6 m1_354_22513# m1_354_22513# m1_31535_22102# m1_31535_22102# m1_31771_21430#
+ vss nfet$383
Xnfet$390_7 m1_n7401_15478# m1_n7401_15478# m1_n927_19404# m1_n927_19404# m1_n695_20470#
+ vss nfet$390
Xnfet$369_4 m1_12259_24224# m1_12259_24224# m1_11903_24542# m1_11903_24542# m1_12357_24542#
+ vss nfet$369
Xnfet$389_18 m1_23930_15778# m1_23930_15778# m1_23820_18030# m1_23820_18030# m1_24056_17358#
+ vss nfet$389
Xnfet$381_3 m1_326_24346# m1_326_24346# vss vss m1_n192_24542# vss nfet$381
Xnfet$374_2 m1_12805_21786# vss m1_12935_21590# vss nfet$374
Xnfet$370_75 m1_28371_23922# vss m1_28991_24224# vss nfet$370
Xpfet$352_16 vdd vdd m1_29256_21786# m1_28624_21786# pfet$352
Xnfet$370_64 m1_19644_25858# vss m1_19781_25662# vss nfet$370
Xnfet$370_53 m1_23827_25858# m1_24451_25662# m1_24188_23922# vss nfet$370
Xnfet$370_42 m1_15943_25858# vss m1_16085_25662# vss nfet$370
Xnfet$370_31 m1_15943_25858# vss m1_18339_24542# vss nfet$370
Xpfet$359_2 vdd m1_30256_19792# vdd m1_24973_22513# pfet$359
Xnfet$370_20 pd3 vss m1_5771_21786# vss nfet$370
Xpfet$366_3 vdd m1_n5461_18030# vdd m1_n6788_16080# pfet$366
Xpfet$373_4 vdd vdd m1_n4485_21904# m1_n3822_21786# pfet$373
Xpfet$364_0 vdd vdd fout m1_34093_22102# pfet$364
Xpfet$352_9 vdd vdd m1_22222_21786# m1_21590_21786# pfet$352
Xpfet$371_1 vdd vdd m1_n6111_25858# m1_n6856_24542# pfet$371
Xpfet$350_6 vdd vdd vdd m1_10505_22402# m1_9288_21786# m1_9288_21786# pfet$350
Xpfet$348_106 vdd vdd m1_25107_21786# m1_28492_25858# pfet$348
Xpfet$348_92 vdd vdd m1_28492_25858# m1_29607_24346# pfet$348
Xpfet$348_81 vdd vdd m1_18339_24542# m1_15943_25858# pfet$348
Xpfet$348_70 vdd vdd m1_14156_24542# m1_11760_25858# pfet$348
Xnfet$399_4 m1_n4623_25487# m1_n2567_23922# m1_n3184_24224# vss nfet$399
Xnfet$378_9 m1_n7513_20152# vss m1_33790_24346# vss nfet$378
Xnfet$373_75 sd3 vss m1_17697_15478# vss nfet$373
Xnfet$373_64 m1_13668_17714# vss m1_13198_17714# vss nfet$373
Xnfet$373_53 m1_22848_17343# vss m1_23007_17836# vss nfet$373
Xnfet$373_31 m1_1933_17343# m1_3989_15778# m1_3372_16080# vss nfet$373
Xnfet$373_20 m1_1119_17714# vss m1_1709_17518# vss nfet$373
Xnfet$373_42 m1_n811_16080# vss m1_n1168_15778# vss nfet$373
Xnfet$397_1 m1_n8625_26174# vss m1_n7082_23622# vss nfet$397
Xnfet$383_7 m1_3871_22513# m1_3871_22513# vss vss m1_31771_21430# vss nfet$383
Xnfet$390_8 m1_26063_15478# m1_26063_15478# m1_n3822_20130# m1_n3822_20130# m1_27441_20470#
+ vss nfet$390
Xnfet$369_5 m1_8692_24346# m1_8692_24346# vss vss m1_8174_24542# vss nfet$369
Xnfet$381_4 m1_33174_24224# m1_33174_24224# m1_32818_24542# m1_32818_24542# m1_33272_24542#
+ vss nfet$381
Xnfet$389_19 m1_23109_16202# m1_23109_16202# vss vss m1_22591_16398# vss nfet$389
Xnfet$374_3 m1_9288_21786# vss m1_9418_21590# vss nfet$374
Xpfet$352_17 vdd vdd m1_25739_21786# m1_25107_21786# pfet$352
Xnfet$370_76 m1_28492_25858# vss m1_28634_25662# vss nfet$370
Xnfet$370_65 m1_28492_25858# vss m1_25107_21786# vss nfet$370
Xnfet$370_54 m1_24309_25858# vss m1_24451_25662# vss nfet$370
Xnfet$370_43 m1_15461_25858# vss m1_15598_25662# vss nfet$370
Xnfet$370_32 m1_15461_25858# m1_17546_25658# m1_18339_24542# vss nfet$370
Xpfet$359_3 vdd vdd m1_34843_21786# m1_34093_19792# pfet$359
Xpfet$366_4 vdd vdd m1_26217_17714# m1_26676_16080# pfet$366
Xnfet$370_21 m1_11278_25858# m1_11902_25662# m1_11639_23922# vss nfet$370
Xnfet$370_10 m1_7577_25858# vss m1_9973_24542# vss nfet$370
Xpfet$373_5 vdd m1_n6839_21786# vdd m1_n5764_21786# pfet$373
Xnfet$372_0 m1_n3534_17714# m1_n3534_17714# vss vss m1_3454_20470# vss nfet$372
Xpfet$357_0 vdd vdd m1_n646_24542# m1_n290_24224# pfet$357
Xpfet$350_7 vdd m1_354_22513# m1_354_22513# m1_n674_22102# m1_1120_21786# m1_1120_21786#
+ pfet$350
Xpfet$348_107 vdd m1_24309_25858# vdd m1_25912_25658# pfet$348
Xpfet$348_93 vdd m1_28991_24224# m1_30095_25658# m1_28010_25858# pfet$348
Xpfet$348_82 vdd vdd m1_21241_24346# m1_n7513_20152# pfet$348
Xpfet$348_71 vdd vdd m1_11039_21786# m1_11760_25858# pfet$348
Xpfet$348_60 vdd vdd m1_20126_25858# m1_21241_24346# pfet$348
Xnfet$399_5 m1_n4464_25980# m1_n3541_23922# m1_n4362_24346# vss nfet$399
Xnfet$373_76 m1_14482_17343# m1_16538_15778# m1_15921_16080# vss nfet$373
Xnfet$373_65 m1_14482_17343# m1_14743_16202# m1_14258_17518# vss nfet$373
Xnfet$373_54 m1_22848_17343# m1_23109_16202# m1_22624_17518# vss nfet$373
Xnfet$373_32 m1_2092_17836# m1_3015_15778# m1_2194_16202# vss nfet$373
Xnfet$373_21 m1_1933_17343# m1_2194_16202# m1_1709_17518# vss nfet$373
Xnfet$373_10 m1_11738_16080# vss m1_11381_15778# vss nfet$373
Xnfet$373_43 sd8 vss m1_n3218_15478# vss nfet$373
Xnfet$397_2 vss vss m1_n9336_24346# vss nfet$397
Xnfet$390_9 m1_29239_20152# m1_29239_20152# m1_n3822_20130# m1_n3822_20130# m1_28073_20470#
+ vss nfet$390
Xnfet$369_6 m1_8076_24224# m1_8076_24224# m1_7720_24542# m1_7720_24542# m1_8174_24542#
+ vss nfet$369
Xnfet$381_5 m1_33790_24346# m1_33790_24346# vss vss m1_33272_24542# vss nfet$381
Xnfet$374_4 m1_7522_21786# vss m1_8154_21786# vss nfet$374
Xnfet$370_77 m1_28010_25858# vss m1_28147_25662# vss nfet$370
Xnfet$370_66 m1_28010_25858# m1_30095_25658# m1_30888_24542# vss nfet$370
Xnfet$370_55 m1_23827_25858# vss m1_23964_25662# vss nfet$370
Xnfet$370_44 m1_15822_23922# vss m1_16442_24224# vss nfet$370
Xnfet$370_33 m1_11760_25858# vss m1_14156_24542# vss nfet$370
Xpfet$359_4 vdd m1_34093_19792# vdd m1_32818_20470# pfet$359
Xpfet$366_5 vdd m1_26217_17714# vdd m1_27292_16202# pfet$366
Xnfet$370_22 m1_11760_25858# vss m1_11902_25662# vss nfet$370
Xnfet$370_11 m1_7522_21786# vss m1_11278_25858# vss nfet$370
Xpfet$373_6 vdd vdd m1_n6973_21481# m1_n6839_21786# pfet$373
Xnfet$372_1 m1_2384_19550# m1_2384_19550# vss vss m1_2822_20470# vss nfet$372
Xpfet$357_1 vdd m1_n789_25858# vdd m1_814_25658# pfet$357
Xpfet$348_108 vdd vdd m1_25424_24346# m1_n7513_20152# pfet$348
Xpfet$350_8 vdd vdd vdd m1_6360_22102# m1_5901_21590# m1_5901_21590# pfet$350
Xpfet$348_94 vdd m1_28492_25858# vdd m1_30095_25658# pfet$348
Xpfet$348_83 vdd m1_21729_25658# m1_22522_24542# m1_19781_25662# pfet$348
Xpfet$348_72 vdd m1_13363_25658# m1_14156_24542# m1_11415_25662# pfet$348
Xpfet$348_61 vdd m1_24452_24542# vdd m1_25424_24346# pfet$348
Xpfet$348_50 vdd vdd m1_20268_25662# m1_20126_25858# pfet$348
Xnfet$399_6 m1_n4464_25980# m1_n3184_24224# m1_n3651_26174# vss nfet$399
Xnfet$397_3 fin vss m1_n10933_25858# vss nfet$397
Xnfet$373_77 sd4 vss m1_13514_15478# vss nfet$373
Xnfet$373_66 m1_n7513_20152# vss m1_14127_16080# vss nfet$373
Xnfet$373_55 m1_22034_17714# vss m1_24904_15778# vss nfet$373
Xnfet$373_44 m1_n2091_17836# m1_n811_16080# m1_n1278_18030# vss nfet$373
Xnfet$373_33 sd7 vss m1_965_15478# vss nfet$373
Xnfet$373_22 m1_6116_17343# m1_6377_16202# m1_5892_17518# vss nfet$373
Xnfet$373_11 m1_10299_17343# m1_12355_15778# m1_11738_16080# vss nfet$373
Xnfet$369_7 m1_9180_25658# m1_9180_25658# vss vss m1_9639_25502# vss nfet$369
Xnfet$395_0 m1_n7082_23622# m1_n6856_24542# vss vss nfet$395
Xnfet$381_6 m1_33790_24346# m1_33790_24346# m1_32675_25947# m1_32675_25947# m1_34737_25502#
+ vss nfet$381
Xnfet$370_78 m1_28010_25858# m1_28634_25662# m1_28371_23922# vss nfet$370
Xnfet$370_67 m1_28492_25858# vss m1_30888_24542# vss nfet$370
Xnfet$370_56 m1_19781_25662# m1_20625_24224# m1_21729_25658# vss nfet$370
Xnfet$370_45 m1_15461_25858# m1_16085_25662# m1_15822_23922# vss nfet$370
Xnfet$370_34 m1_11278_25858# m1_13363_25658# m1_14156_24542# vss nfet$370
Xpfet$366_6 vdd vdd m1_28003_18030# m1_28113_15778# pfet$366
Xpfet$359_5 vdd vdd m1_34093_19792# m1_32818_21586# pfet$359
Xnfet$370_23 m1_11278_25858# vss m1_11415_25662# vss nfet$370
Xnfet$370_12 m1_7577_25858# vss m1_7522_21786# vss nfet$370
Xpfet$373_7 vdd vdd m1_n6839_21786# m1_n6380_21786# pfet$373
Xnfet$374_5 m1_488_21786# vss m1_1120_21786# vss nfet$374
Xnfet$372_2 m1_5901_19550# m1_5901_19550# vss vss m1_6339_20470# vss nfet$372
Xpfet$357_2 vdd vdd m1_n789_25858# m1_326_24346# pfet$357
Xpfet$348_109 vdd m1_12259_24224# m1_13363_25658# m1_11278_25858# pfet$348
Xpfet$350_9 vdd m1_3871_22513# m1_3871_22513# m1_3471_22402# m1_4005_21786# m1_4005_21786#
+ pfet$350
Xpfet$362_0 vdd m1_34093_22102# vdd m1_28490_22513# pfet$362
Xnfet$399_7 m1_n4623_25487# m1_n4362_24346# m1_n4847_25662# vss nfet$399
Xpfet$348_95 vdd vdd m1_28991_24224# m1_28371_23922# pfet$348
Xpfet$348_84 vdd vdd m1_23827_25858# m1_18073_21786# pfet$348
Xpfet$348_73 vdd m1_16086_24542# vdd m1_17058_24346# pfet$348
Xpfet$348_62 vdd vdd m1_24452_24542# m1_24808_24224# pfet$348
Xpfet$348_51 vdd vdd m1_20625_24224# m1_20005_23922# pfet$348
Xpfet$348_40 vdd vdd m1_11760_25858# m1_12875_24346# pfet$348
Xpfet$350_30 vdd vdd vdd m1_17539_22402# m1_16322_21786# m1_16322_21786# pfet$350
Xnfet$397_4 m1_n10572_23922# vss m1_n9952_24224# vss nfet$397
Xnfet$373_78 m1_14641_17836# m1_15564_15778# m1_14743_16202# vss nfet$373
Xnfet$373_67 m1_17381_17714# vss m1_14482_17343# vss nfet$373
Xnfet$373_56 m1_24287_16080# vss m1_23930_15778# vss nfet$373
Xnfet$373_45 m1_n3064_17714# vss m1_n194_15778# vss nfet$373
Xnfet$373_34 m1_n2250_17343# vss m1_n2091_17836# vss nfet$373
Xnfet$373_23 m1_5302_17714# vss m1_4832_17714# vss nfet$373
Xnfet$373_12 m1_9485_17714# vss m1_12355_15778# vss nfet$373
Xnfet$369_8 m1_8692_24346# m1_8692_24346# m1_7577_25858# m1_7577_25858# m1_9639_25502#
+ vss nfet$369
Xnfet$388_0 fout vss m1_35837_22102# vss nfet$388
Xnfet$395_1 m1_n8283_19850# vss m1_n6856_24542# vss nfet$395
Xnfet$381_7 m1_34278_25658# m1_34278_25658# vss vss m1_34737_25502# vss nfet$381
Xnfet$370_57 m1_20126_25858# vss m1_20268_25662# vss nfet$370
Xnfet$370_46 m1_20126_25858# vss m1_18073_21786# vss nfet$370
Xnfet$370_35 m1_15598_25662# m1_15822_23922# m1_16086_24542# vss nfet$370
Xpfet$366_7 vdd m1_28003_18030# vdd m1_26676_16080# pfet$366
Xnfet$370_24 m1_7095_25858# m1_7719_25662# m1_7456_23922# vss nfet$370
Xnfet$370_13 m1_11415_25662# m1_11639_23922# m1_11903_24542# vss nfet$370
Xnfet$374_6 m1_5771_21786# vss m1_5901_21590# vss nfet$374
Xnfet$370_79 pd7 vss m1_19839_21786# vss nfet$370
Xnfet$370_68 m1_n7513_20152# vss m1_29607_24346# vss nfet$370
Xpfet$359_6 vdd vdd m1_31535_19792# m1_14422_22513# pfet$359
Xnfet$372_3 m1_4832_17714# m1_4832_17714# vss vss m1_10488_20470# vss nfet$372
Xpfet$357_3 vdd m1_n646_24542# vdd m1_326_24346# pfet$357
Xnfet$370_0 m1_3394_25858# vss m1_5790_24542# vss nfet$370
Xpfet$362_1 vdd vdd m1_34093_22102# m1_34843_21786# pfet$362
Xpfet$355_0 vdd vdd m1_n7401_15478# sd9 pfet$355
Xpfet$348_96 vdd m1_28635_24542# vdd m1_29607_24346# pfet$348
Xpfet$348_85 vdd m1_24188_23922# m1_24452_24542# m1_23827_25858# pfet$348
Xpfet$348_74 vdd vdd m1_14556_21786# m1_15943_25858# pfet$348
Xpfet$348_63 vdd vdd m1_19781_25662# m1_19644_25858# pfet$348
Xpfet$348_52 vdd m1_20268_25662# m1_20005_23922# m1_19781_25662# pfet$348
Xpfet$348_41 vdd vdd m1_9288_21786# pd4 pfet$348
Xpfet$348_30 vdd vdd m1_2912_25858# m1_488_21786# pfet$348
Xpfet$350_31 vdd vdd vdd m1_27462_22102# m1_27003_21590# m1_27003_21590# pfet$350
Xpfet$350_20 vdd vdd vdd m1_20428_22102# m1_19969_21590# m1_19969_21590# pfet$350
Xnfet$397_5 m1_n10933_25858# vss m1_n10796_25662# vss nfet$397
Xnfet$373_79 m1_15921_16080# vss m1_15564_15778# vss nfet$373
Xnfet$373_68 m1_18665_17343# m1_18926_16202# m1_18441_17518# vss nfet$373
Xnfet$373_57 m1_22848_17343# m1_24904_15778# m1_24287_16080# vss nfet$373
Xnfet$373_46 m1_22034_17714# vss m1_21564_17714# vss nfet$373
Xnfet$373_24 m1_4832_17714# vss m1_1933_17343# vss nfet$373
Xnfet$373_13 m1_10458_17836# m1_11381_15778# m1_10560_16202# vss nfet$373
Xnfet$373_35 m1_n7513_20152# vss m1_5761_16080# vss nfet$373
Xnfet$369_9 m1_17058_24346# m1_17058_24346# vss vss m1_16540_24542# vss nfet$369
Xnfet$388_1 define m1_35837_22102# vss vss nfet$388
Xnfet$374_7 m1_4005_21786# vss m1_4637_21786# vss nfet$374
Xpfet$359_7 vdd vdd m1_31535_22102# m1_354_22513# pfet$359
Xnfet$370_69 m1_24309_25858# vss m1_26705_24542# vss nfet$370
Xnfet$370_58 m1_20005_23922# vss m1_20625_24224# vss nfet$370
Xnfet$370_47 m1_23964_25662# m1_24188_23922# m1_24452_24542# vss nfet$370
Xnfet$370_36 m1_11760_25858# vss m1_11039_21786# vss nfet$370
Xnfet$370_25 m1_7232_25662# m1_8076_24224# m1_9180_25658# vss nfet$370
Xnfet$370_14 m1_n7513_20152# vss m1_8692_24346# vss nfet$370
Xpfet$357_4 vdd vdd m1_32675_25947# m1_33790_24346# pfet$357
Xnfet$372_4 m1_9418_19550# m1_9418_19550# vss vss m1_9856_20470# vss nfet$372
Xnfet$370_1 m1_2912_25858# m1_4997_25658# m1_5790_24542# vss nfet$370
Xpfet$362_2 vdd vdd m1_30256_22102# m1_7388_22513# pfet$362
Xpfet$355_1 vdd vdd m1_21880_15478# sd2 pfet$355
Xpfet$348_0 vdd vdd m1_3049_25662# m1_2912_25858# pfet$348
Xpfet$348_97 vdd vdd m1_21590_21786# m1_24309_25858# pfet$348
Xpfet$348_86 vdd m1_28634_25662# m1_28371_23922# m1_28147_25662# pfet$348
Xpfet$348_75 vdd vdd m1_19644_25858# m1_14556_21786# pfet$348
Xpfet$348_64 vdd vdd m1_22522_24542# m1_20126_25858# pfet$348
Xpfet$348_53 vdd m1_20625_24224# m1_21729_25658# m1_19644_25858# pfet$348
Xpfet$348_42 vdd m1_11760_25858# vdd m1_13363_25658# pfet$348
Xpfet$348_31 vdd m1_3273_23922# m1_3537_24542# m1_2912_25858# pfet$348
Xpfet$348_20 vdd vdd m1_4509_24346# m1_n7513_20152# pfet$348
Xpfet$350_32 vdd m1_28490_22513# m1_28490_22513# m1_28090_22402# m1_28624_21786# m1_28624_21786#
+ pfet$350
Xpfet$350_21 vdd vdd vdd m1_21056_22402# m1_19839_21786# m1_19839_21786# pfet$350
Xpfet$350_10 vdd m1_3871_22513# m1_3871_22513# m1_2843_22102# m1_4637_21786# m1_4637_21786#
+ pfet$350
Xnfet$373_69 m1_17851_17714# vss m1_17381_17714# vss nfet$373
Xnfet$373_58 m1_23007_17836# m1_23930_15778# m1_23109_16202# vss nfet$373
Xnfet$373_47 m1_22034_17714# vss m1_22624_17518# vss nfet$373
Xnfet$373_25 m1_2092_17836# m1_3372_16080# m1_2905_18030# vss nfet$373
Xnfet$373_14 m1_6116_17343# m1_8172_15778# m1_7555_16080# vss nfet$373
Xnfet$373_36 m1_n3064_17714# vss m1_n2474_17518# vss nfet$373
Xnfet$397_6 m1_n10452_25858# vss m1_n10309_25662# vss nfet$397
Xnfet$374_8 m1_2254_21786# vss m1_2384_21590# vss nfet$374
Xnfet$370_59 m1_19644_25858# m1_20268_25662# m1_20005_23922# vss nfet$370
Xnfet$370_48 m1_18073_21786# vss m1_23827_25858# vss nfet$370
Xnfet$370_37 m1_11039_21786# vss m1_15461_25858# vss nfet$370
Xnfet$370_26 m1_7095_25858# m1_9180_25658# m1_9973_24542# vss nfet$370
Xnfet$370_15 m1_7232_25662# m1_7456_23922# m1_7720_24542# vss nfet$370
Xnfet$393_0 m1_n5351_15778# m1_n5351_15778# m1_n5461_18030# m1_n5461_18030# m1_n5225_17358#
+ vss nfet$393
Xpfet$378_0 vdd vdd m1_n5227_20152# m1_n2543_20130# pfet$378
Xnfet$372_5 m1_649_17714# m1_649_17714# vss vss m1_6971_20470# vss nfet$372
Xpfet$357_5 vdd m1_32675_25947# vdd m1_34278_25658# pfet$357
Xpfet$353_10 vdd vdd m1_27031_17343# m1_n10452_25858# pfet$353
Xnfet$370_2 m1_n7513_20152# vss m1_4509_24346# vss nfet$370
Xpfet$355_2 vdd vdd m1_26063_15478# sd1 pfet$355
Xpfet$362_3 vdd m1_31535_22102# vdd m1_3871_22513# pfet$362
Xpfet$348_1 vdd m1_3536_25662# m1_3273_23922# m1_3049_25662# pfet$348
Xpfet$348_98 vdd m1_30095_25658# m1_30888_24542# m1_28147_25662# pfet$348
Xpfet$348_87 vdd vdd m1_28147_25662# m1_28010_25858# pfet$348
Xpfet$348_76 vdd m1_20005_23922# m1_20269_24542# m1_19644_25858# pfet$348
Xpfet$348_65 vdd vdd m1_18073_21786# m1_20126_25858# pfet$348
Xpfet$348_54 vdd vdd m1_24808_24224# m1_24188_23922# pfet$348
Xpfet$348_43 vdd vdd m1_12805_21786# pd5 pfet$348
Xpfet$348_32 vdd vdd m1_7720_24542# m1_8076_24224# pfet$348
Xpfet$348_21 vdd m1_7456_23922# m1_7720_24542# m1_7095_25858# pfet$348
Xpfet$348_10 vdd m1_8076_24224# m1_9180_25658# m1_7095_25858# pfet$348
Xpfet$350_33 vdd m1_28490_22513# m1_28490_22513# m1_27462_22102# m1_29256_21786# m1_29256_21786#
+ pfet$350
Xpfet$350_22 vdd m1_21456_22513# m1_21456_22513# m1_20428_22102# m1_22222_21786# m1_22222_21786#
+ pfet$350
Xpfet$360_0 vdd m1_n647_25662# m1_n910_23922# m1_n1134_25662# pfet$360
Xpfet$350_11 vdd vdd vdd m1_2843_22102# m1_2384_21590# m1_2384_21590# pfet$350
Xnfet$373_59 m1_17851_17714# vss m1_20721_15778# vss nfet$373
Xnfet$373_48 m1_18824_17836# m1_20104_16080# m1_19637_18030# vss nfet$373
Xnfet$373_26 m1_5302_17714# vss m1_5892_17518# vss nfet$373
Xnfet$373_15 m1_5302_17714# vss m1_8172_15778# vss nfet$373
Xnfet$373_37 m1_n7513_20152# vss m1_n2605_16080# vss nfet$373
Xnfet$397_7 m1_n7320_25516# vss m1_n2567_23922# vss nfet$397
Xpfet$356_10 vdd vdd m1_35071_24542# m1_32675_25947# pfet$356
Xnfet$374_9 m1_23356_21786# vss m1_23486_21590# vss nfet$374
Xnfet$370_49 m1_19781_25662# m1_20005_23922# m1_20269_24542# vss nfet$370
Xnfet$370_38 m1_n7513_20152# vss m1_12875_24346# vss nfet$370
Xnfet$386_0 m1_34093_19792# vss m1_34843_21786# vss nfet$386
Xnfet$370_27 m1_7577_25858# vss m1_7719_25662# vss nfet$370
Xnfet$370_16 m1_4005_21786# vss m1_7095_25858# vss nfet$370
Xnfet$393_1 m1_n6788_16080# m1_n6788_16080# vss vss m1_n5225_17358# vss nfet$393
Xpfet$378_1 vdd m1_n4485_20152# vdd m1_n3206_20274# pfet$378
Xnfet$372_6 m1_n1133_19550# m1_n1133_19550# vss vss m1_n695_20470# vss nfet$372
Xpfet$357_6 vdd vdd m1_32818_24542# m1_33174_24224# pfet$357
Xpfet$353_11 vdd vdd m1_26807_17518# m1_26217_17714# pfet$353
Xpfet$362_4 vdd m1_30256_22102# vdd m1_9645_21447# pfet$362
Xnfet$370_3 m1_488_21786# vss m1_2912_25858# vss nfet$370
Xpfet$348_99 vdd vdd m1_26705_24542# m1_24309_25858# pfet$348
Xpfet$348_88 vdd vdd m1_28634_25662# m1_28492_25858# pfet$348
Xpfet$348_77 vdd vdd m1_20269_24542# m1_20625_24224# pfet$348
Xpfet$348_66 vdd vdd m1_15461_25858# m1_11039_21786# pfet$348
Xpfet$348_55 vdd m1_24451_25662# m1_24188_23922# m1_23964_25662# pfet$348
Xpfet$348_44 vdd m1_15943_25858# vdd m1_17546_25658# pfet$348
Xpfet$348_33 vdd vdd m1_7522_21786# m1_7577_25858# pfet$348
Xpfet$348_22 vdd vdd m1_3537_24542# m1_3893_24224# pfet$348
Xpfet$348_11 vdd vdd m1_7719_25662# m1_7577_25858# pfet$348
Xpfet$348_2 vdd vdd m1_3394_25858# m1_4509_24346# pfet$348
Xpfet$353_0 vdd vdd m1_n6274_17836# m1_n6433_17343# pfet$353
Xpfet$360_1 vdd m1_n910_23922# m1_n646_24542# m1_n1271_25858# pfet$360
Xpfet$350_34 vdd vdd vdd m1_28090_22402# m1_26873_21786# m1_26873_21786# pfet$350
Xpfet$350_23 vdd vdd vdd m1_23945_22102# m1_23486_21590# m1_23486_21590# pfet$350
Xnfet$397_8 m1_n4623_25487# vss m1_n4464_25980# vss nfet$397
Xpfet$350_12 vdd vdd vdd m1_3471_22402# m1_2254_21786# m1_2254_21786# pfet$350
Xnfet$373_49 m1_21564_17714# vss m1_18665_17343# vss nfet$373
Xnfet$373_27 m1_1119_17714# vss m1_3989_15778# vss nfet$373
Xnfet$373_16 m1_6275_17836# m1_7198_15778# m1_6377_16202# vss nfet$373
Xnfet$373_38 m1_n2250_17343# m1_n1989_16202# m1_n2474_17518# vss nfet$373
Xpfet$356_11 vdd vdd m1_32817_25662# m1_32675_25947# pfet$356
Xnfet$370_39 pd4 vss m1_9288_21786# vss nfet$370
Xnfet$386_1 m1_30256_19792# vss m1_32818_20470# vss nfet$386
Xnfet$370_28 m1_3394_25858# vss m1_4005_21786# vss nfet$370
Xnfet$370_17 m1_11639_23922# vss m1_12259_24224# vss nfet$370
Xnfet$393_2 m1_n6788_16080# m1_n6788_16080# m1_n7247_17714# m1_n7247_17714# m1_n6690_16398#
+ vss nfet$393
Xnfet$379_0 m1_n1134_25662# m1_n910_23922# m1_n646_24542# vss nfet$379
Xpfet$378_2 vdd m1_n5227_20152# vdd m1_n1927_20274# pfet$378
Xnfet$372_7 m1_n7383_17599# m1_n7383_17599# vss vss m1_n63_20470# vss nfet$372
Xpfet$357_7 vdd m1_32818_24542# vdd m1_33790_24346# pfet$357
Xpfet$353_12 vdd vdd m1_26676_16080# m1_n7513_20152# pfet$353
Xnfet$370_4 m1_2912_25858# vss m1_3049_25662# vss nfet$370
Xpfet$348_34 vdd m1_9180_25658# m1_9973_24542# m1_7232_25662# pfet$348
Xpfet$348_23 vdd m1_3537_24542# vdd m1_4509_24346# pfet$348
Xpfet$348_12 vdd m1_7577_25858# vdd m1_9180_25658# pfet$348
Xpfet$348_3 vdd m1_3394_25858# vdd m1_4997_25658# pfet$348
Xpfet$348_89 vdd vdd m1_19839_21786# pd7 pfet$348
Xpfet$348_78 vdd m1_20269_24542# vdd m1_21241_24346# pfet$348
Xpfet$348_67 vdd m1_15822_23922# m1_16086_24542# m1_15461_25858# pfet$348
Xpfet$348_56 vdd m1_24808_24224# m1_25912_25658# m1_23827_25858# pfet$348
Xpfet$348_45 vdd vdd m1_16442_24224# m1_15822_23922# pfet$348
Xpfet$353_1 vdd vdd m1_n4377_15778# m1_n7247_17714# pfet$353
Xpfet$360_2 vdd m1_n290_24224# m1_814_25658# m1_n1271_25858# pfet$360
Xpfet$350_35 vdd vdd vdd m1_13394_22102# m1_12935_21590# m1_12935_21590# pfet$350
Xpfet$350_24 vdd m1_17939_22513# m1_17939_22513# m1_16911_22102# m1_18705_21786# m1_18705_21786#
+ pfet$350
Xpfet$350_13 vdd vdd vdd m1_6988_22402# m1_5771_21786# m1_5771_21786# pfet$350
Xnfet$397_9 m1_n3184_24224# vss m1_n3541_23922# vss nfet$397
Xnfet$373_28 m1_1933_17343# vss m1_2092_17836# vss nfet$373
Xnfet$373_17 m1_649_17714# vss m1_n2250_17343# vss nfet$373
Xnfet$373_39 m1_n3064_17714# vss m1_n3534_17714# vss nfet$373
Xpfet$356_12 vdd vdd m1_32193_25858# m1_25107_21786# pfet$356
Xnfet$370_29 m1_15943_25858# vss m1_14556_21786# vss nfet$370
Xnfet$370_18 m1_7095_25858# vss m1_7232_25662# vss nfet$370
Xnfet$393_3 m1_n6172_16202# m1_n6172_16202# vss vss m1_n6690_16398# vss nfet$393
Xnfet$386_2 m1_31535_19792# m1_32818_20470# vss vss nfet$386
Xpfet$378_3 vdd m1_n6839_20152# vdd m1_n927_19404# pfet$378
Xnfet$379_1 m1_n1271_25858# m1_n647_25662# m1_n910_23922# vss nfet$379
Xnfet$372_8 m1_27003_19550# m1_27003_19550# vss vss m1_27441_20470# vss nfet$372
Xnfet$391_0 m1_35837_22102# vss m1_n7513_20152# vss nfet$391
Xpfet$353_13 vdd vdd m1_25747_17714# m1_26217_17714# pfet$353
Xpfet$376_0 vdd vdd vdd m1_n8047_19550# m1_n7513_20152# m1_n7513_20152# pfet$376
Xnfet$370_5 m1_2912_25858# m1_3536_25662# m1_3273_23922# vss nfet$370
Xpfet$348_4 vdd vdd m1_3893_24224# m1_3273_23922# pfet$348
Xnfet$404_0 m1_n4485_20152# m1_n6380_21786# vss vss nfet$404
Xpfet$348_79 vdd m1_17546_25658# m1_18339_24542# m1_15598_25662# pfet$348
Xpfet$348_68 vdd vdd m1_16086_24542# m1_16442_24224# pfet$348
Xpfet$348_57 vdd vdd m1_24451_25662# m1_24309_25858# pfet$348
Xpfet$348_46 vdd m1_16442_24224# m1_17546_25658# m1_15461_25858# pfet$348
Xpfet$348_35 vdd m1_7720_24542# vdd m1_8692_24346# pfet$348
Xpfet$348_24 vdd vdd m1_5790_24542# m1_3394_25858# pfet$348
Xpfet$348_13 vdd vdd m1_12259_24224# m1_11639_23922# pfet$348
Xpfet$360_3 vdd m1_814_25658# m1_1607_24542# m1_n1134_25662# pfet$360
Xpfet$353_2 vdd vdd m1_n5351_15778# m1_n4994_16080# pfet$353
Xpfet$350_25 vdd m1_17939_22513# m1_17939_22513# m1_17539_22402# m1_18073_21786# m1_18073_21786#
+ pfet$350
Xpfet$350_14 vdd vdd vdd m1_n46_22402# m1_n1263_21786# m1_n1263_21786# pfet$350
Xnfet$373_29 m1_3372_16080# vss m1_3015_15778# vss nfet$373
Xnfet$373_18 m1_1119_17714# vss m1_649_17714# vss nfet$373
Xpfet$356_13 vdd vdd m1_33790_24346# m1_n7513_20152# pfet$356
Xnfet$386_3 m1_30256_22102# vss m1_32818_21586# vss nfet$386
Xnfet$393_4 m1_28113_15778# m1_28113_15778# m1_28003_18030# m1_28003_18030# m1_28239_17358#
+ vss nfet$393
Xnfet$370_19 m1_7456_23922# vss m1_8076_24224# vss nfet$370
Xpfet$378_4 vdd vdd m1_n6839_20152# m1_n6973_21481# pfet$378
Xnfet$379_2 m1_n1271_25858# m1_814_25658# m1_1607_24542# vss nfet$379
Xnfet$384_0 m1_34843_21786# m1_34843_21786# m1_34093_22102# m1_34093_22102# m1_34329_21430#
+ vss nfet$384
Xnfet$372_9 m1_25747_17714# m1_25747_17714# vss vss m1_28073_20470# vss nfet$372
Xpfet$376_1 vdd m1_n8283_19850# m1_n8283_19850# m1_n8047_19550# m1_n8283_20611# m1_n8283_20611#
+ pfet$376
Xpfet$369_0 vdd vdd vdd m1_n6624_23622# m1_n7082_23622# m1_n7082_23622# pfet$369
Xnfet$370_6 m1_3049_25662# m1_3893_24224# m1_4997_25658# vss nfet$370
Xpfet$348_5 vdd m1_3893_24224# m1_4997_25658# m1_2912_25858# pfet$348
Xnfet$404_1 m1_n5227_20152# vss m1_n6380_21786# vss nfet$404
Xpfet$348_69 vdd vdd m1_12875_24346# m1_n7513_20152# pfet$348
Xpfet$348_58 vdd vdd m1_23964_25662# m1_23827_25858# pfet$348
Xpfet$348_47 vdd vdd m1_15943_25858# m1_17058_24346# pfet$348
Xpfet$348_36 vdd vdd m1_8692_24346# m1_n7513_20152# pfet$348
Xpfet$348_25 vdd vdd m1_4005_21786# m1_3394_25858# pfet$348
Xpfet$348_14 vdd vdd m1_11902_25662# m1_11760_25858# pfet$348
Xpfet$360_4 vdd m1_33174_24224# m1_34278_25658# m1_32193_25858# pfet$360
Xpfet$350_26 vdd vdd vdd m1_16911_22102# m1_16452_21590# m1_16452_21590# pfet$350
Xpfet$350_15 vdd m1_354_22513# m1_354_22513# m1_n46_22402# m1_488_21786# m1_488_21786#
+ pfet$350
Xpfet$353_3 vdd vdd m1_n6657_17518# m1_n7247_17714# pfet$353
Xpfet$349_90 vdd m1_19747_15778# m1_18926_16202# m1_18665_17343# pfet$349
Xnfet$373_19 m1_n7513_20152# vss m1_1578_16080# vss nfet$373
Xpfet$351_0 vdd m1_2590_19404# m1_2590_19404# m1_3458_19550# m1_n3534_17714# m1_n3534_17714#
+ pfet$351
Xnfet$393_5 m1_26676_16080# m1_26676_16080# vss vss m1_28239_17358# vss nfet$393
Xnfet$379_3 m1_n1134_25662# m1_n290_24224# m1_814_25658# vss nfet$379
Xnfet$384_1 m1_28490_22513# m1_28490_22513# vss vss m1_34329_21430# vss nfet$384
Xnfet$377_0 m1_n3534_17714# vss m1_n6433_17343# vss nfet$377
Xpfet$376_2 vdd m1_n8283_20611# m1_n8283_20611# m1_n8047_22344# m1_n8145_21908# m1_n8145_21908#
+ pfet$376
Xpfet$369_1 vdd m1_n6856_24542# m1_n6856_24542# m1_n6624_23622# m1_n8283_19850# m1_n8283_19850#
+ pfet$369
Xnfet$370_7 m1_3049_25662# m1_3273_23922# m1_3537_24542# vss nfet$370
Xpfet$348_6 vdd vdd m1_3536_25662# m1_3394_25858# pfet$348
Xpfet$348_59 vdd vdd m1_16322_21786# pd6 pfet$348
Xpfet$348_48 vdd m1_16085_25662# m1_15822_23922# m1_15598_25662# pfet$348
Xpfet$348_37 vdd vdd m1_9973_24542# m1_7577_25858# pfet$348
Xpfet$348_26 vdd m1_4997_25658# m1_5790_24542# m1_3049_25662# pfet$348
Xpfet$348_15 vdd m1_11902_25662# m1_11639_23922# m1_11415_25662# pfet$348
Xpfet$360_5 vdd m1_32817_25662# m1_32554_23922# m1_32330_25662# pfet$360
Xpfet$350_27 vdd m1_14422_22513# m1_14422_22513# m1_14022_22402# m1_14556_21786# m1_14556_21786#
+ pfet$350
Xpfet$350_16 vdd m1_24973_22513# m1_24973_22513# m1_23945_22102# m1_25739_21786# m1_25739_21786#
+ pfet$350
Xpfet$353_4 vdd vdd m1_n6433_17343# m1_n3534_17714# pfet$353
Xpfet$349_91 vdd m1_24287_16080# m1_23820_18030# m1_22848_17343# pfet$349
Xpfet$349_80 vdd vdd m1_15564_15778# m1_15921_16080# pfet$349
Xpfet$351_1 vdd vdd vdd m1_2822_19850# m1_4620_20152# m1_4620_20152# pfet$351
Xnfet$379_4 m1_32193_25858# m1_34278_25658# m1_35071_24542# vss nfet$379
Xnfet$393_6 m1_27292_16202# m1_27292_16202# vss vss m1_26774_16398# vss nfet$393
Xnfet$384_2 m1_9645_21447# m1_9645_21447# vss vss m1_30492_21430# vss nfet$384
Xnfet$377_1 m1_n7513_20152# vss m1_n6788_16080# vss nfet$377
Xpfet$376_3 vdd vdd vdd m1_n8047_22344# m1_n8283_19850# m1_n8283_19850# pfet$376
Xpfet$348_7 vdd vdd m1_7232_25662# m1_7095_25858# pfet$348
Xnfet$370_8 m1_3394_25858# vss m1_3536_25662# vss nfet$370
Xpfet$348_49 vdd m1_20126_25858# vdd m1_21729_25658# pfet$348
Xpfet$348_38 vdd vdd m1_16085_25662# m1_15943_25858# pfet$348
Xpfet$348_27 vdd vdd m1_11278_25858# m1_7522_21786# pfet$348
Xpfet$348_16 vdd vdd m1_5771_21786# pd3 pfet$348
Xpfet$374_0 vdd vdd m1_n10796_25662# m1_n10933_25858# pfet$374
Xpfet$360_6 vdd m1_34278_25658# m1_35071_24542# m1_32330_25662# pfet$360
Xpfet$353_5 vdd vdd m1_n6788_16080# m1_n7513_20152# pfet$353
Xnfet$402_0 m1_n4485_21904# m1_n5764_21786# vss vss nfet$402
Xpfet$350_28 vdd m1_14422_22513# m1_14422_22513# m1_13394_22102# m1_15188_21786# m1_15188_21786#
+ pfet$350
Xpfet$350_17 vdd m1_21456_22513# m1_21456_22513# m1_21056_22402# m1_21590_21786# m1_21590_21786#
+ pfet$350
Xpfet$349_92 vdd m1_15454_18030# vdd m1_14127_16080# pfet$349
Xpfet$349_81 vdd vdd m1_13668_17714# m1_14127_16080# pfet$349
Xpfet$349_70 vdd vdd m1_18824_17836# m1_18665_17343# pfet$349
Xpfet$351_2 vdd m1_2590_19404# m1_2590_19404# m1_2822_19850# m1_2384_19550# m1_2384_19550#
+ pfet$351
Xnfet$379_5 m1_32330_25662# m1_33174_24224# m1_34278_25658# vss nfet$379
Xnfet$393_7 m1_26676_16080# m1_26676_16080# m1_26217_17714# m1_26217_17714# m1_26774_16398#
+ vss nfet$393
Xnfet$369_20 m1_21241_24346# m1_21241_24346# m1_20126_25858# m1_20126_25858# m1_22188_25502#
+ vss nfet$369
Xnfet$384_3 m1_7388_22513# m1_7388_22513# m1_30256_22102# m1_30256_22102# m1_30492_21430#
+ vss nfet$384
Xnfet$377_2 m1_n4994_16080# vss m1_n5351_15778# vss nfet$377
Xnfet$371_10 m1_19839_21786# m1_19839_21786# m1_21456_22513# m1_21456_22513# m1_21060_21586#
+ vss nfet$371
Xnfet$370_9 m1_3273_23922# vss m1_3893_24224# vss nfet$370
Xpfet$348_39 vdd vdd m1_15598_25662# m1_15461_25858# pfet$348
Xpfet$348_28 vdd m1_11639_23922# m1_11903_24542# m1_11278_25858# pfet$348
Xpfet$348_17 vdd vdd m1_7577_25858# m1_8692_24346# pfet$348
Xpfet$348_8 vdd vdd m1_8076_24224# m1_7456_23922# pfet$348
Xpfet$367_0 vdd m1_n4377_15778# m1_n4994_16080# m1_n6274_17836# pfet$367
Xpfet$374_1 vdd vdd m1_n10309_25662# m1_n10452_25858# pfet$374
Xnfet$382_0 m1_11039_21786# m1_11039_21786# vss vss m1_9877_21586# vss nfet$382
Xpfet$360_7 vdd m1_32554_23922# m1_32818_24542# m1_32193_25858# pfet$360
Xpfet$353_6 vdd vdd m1_n7383_17599# m1_n7247_17714# pfet$353
Xnfet$402_1 m1_n5227_21418# vss m1_n5764_21786# vss nfet$402
Xpfet$350_29 vdd vdd vdd m1_14022_22402# m1_12805_21786# m1_12805_21786# pfet$350
Xpfet$350_18 vdd vdd vdd m1_24573_22402# m1_23356_21786# m1_23356_21786# pfet$350
Xpfet$349_93 vdd m1_23820_18030# vdd m1_22493_16080# pfet$349
Xpfet$349_82 vdd m1_13668_17714# vdd m1_14743_16202# pfet$349
Xpfet$349_71 vdd vdd m1_19747_15778# m1_20104_16080# pfet$349
Xpfet$349_60 vdd vdd m1_n194_15778# m1_n3064_17714# pfet$349
Xpfet$351_3 vdd vdd vdd m1_3458_19550# m1_n3218_15478# m1_n3218_15478# pfet$351
Xnfet$374_10 m1_21590_21786# vss m1_22222_21786# vss nfet$374
Xnfet$379_6 m1_32193_25858# m1_32817_25662# m1_32554_23922# vss nfet$379
Xnfet$369_21 m1_28991_24224# m1_28991_24224# m1_28635_24542# m1_28635_24542# m1_29089_24542#
+ vss nfet$369
Xnfet$369_10 m1_17546_25658# m1_17546_25658# vss vss m1_18005_25502# vss nfet$369
Xnfet$377_3 m1_n6433_17343# vss m1_n6274_17836# vss nfet$377
Xnfet$371_11 m1_19969_21590# m1_19969_21590# m1_21456_22513# m1_21456_22513# m1_20428_21586#
+ vss nfet$371
Xnfet$382_10 m1_21590_21786# m1_21590_21786# vss vss m1_20428_21586# vss nfet$382
Xpfet$348_9 vdd m1_7719_25662# m1_7456_23922# m1_7232_25662# pfet$348
Xnfet$375_0 m1_n3534_17714# vss m1_2384_19550# vss nfet$375
Xnfet$382_1 m1_11671_21786# m1_11671_21786# vss vss m1_10509_21586# vss nfet$382
Xpfet$348_29 vdd vdd m1_11903_24542# m1_12259_24224# pfet$348
Xpfet$348_18 vdd vdd m1_11415_25662# m1_11278_25858# pfet$348
Xpfet$367_1 vdd m1_n5351_15778# m1_n6172_16202# m1_n6433_17343# pfet$367
Xpfet$374_2 vdd vdd m1_n9952_24224# m1_n10572_23922# pfet$374
Xpfet$353_7 vdd vdd m1_27190_17836# m1_27031_17343# pfet$353
Xnfet$402_2 m1_n6839_21786# vss m1_n6973_21481# vss nfet$402
Xpfet$350_19 vdd m1_24973_22513# m1_24973_22513# m1_24573_22402# m1_25107_21786# m1_25107_21786#
+ pfet$350
Xnfet$377_10 m1_26217_17714# vss m1_29087_15778# vss nfet$377
Xpfet$349_94 vdd vdd m1_22624_17518# m1_22034_17714# pfet$349
Xpfet$349_83 vdd m1_16538_15778# m1_15921_16080# m1_14641_17836# pfet$349
Xpfet$349_72 vdd m1_20721_15778# m1_20104_16080# m1_18824_17836# pfet$349
Xpfet$349_61 vdd m1_n811_16080# m1_n1278_18030# m1_n2250_17343# pfet$349
Xpfet$349_50 vdd m1_n1168_15778# m1_n1989_16202# m1_n2250_17343# pfet$349
Xpfet$351_4 vdd m1_6107_19404# m1_6107_19404# m1_6339_19850# m1_5901_19550# m1_5901_19550#
+ pfet$351
Xnfet$374_11 m1_18073_21786# vss m1_18705_21786# vss nfet$374
Xnfet$390_10 m1_9331_15478# m1_9331_15478# m1_n3822_21786# m1_n3822_21786# m1_13373_20470#
+ vss nfet$390
Xnfet$379_7 m1_32330_25662# m1_32554_23922# m1_32818_24542# vss nfet$379
Xnfet$369_22 m1_29607_24346# m1_29607_24346# vss vss m1_29089_24542# vss nfet$369
Xnfet$369_11 m1_16442_24224# m1_16442_24224# m1_16086_24542# m1_16086_24542# m1_16540_24542#
+ vss nfet$369
Xnfet$377_4 m1_n7247_17714# vss m1_n4377_15778# vss nfet$377
Xnfet$371_12 m1_16322_21786# m1_16322_21786# m1_17939_22513# m1_17939_22513# m1_17543_21586#
+ vss nfet$371
Xnfet$375_1 m1_n3218_15478# vss m1_4620_20152# vss nfet$375
Xnfet$382_2 m1_8154_21786# m1_8154_21786# vss vss m1_6992_21586# vss nfet$382
Xnfet$382_11 m1_22222_21786# m1_22222_21786# vss vss m1_21060_21586# vss nfet$382
Xpfet$348_19 vdd vdd m1_7095_25858# m1_4005_21786# pfet$348
Xpfet$367_2 vdd m1_n4994_16080# m1_n5461_18030# m1_n6433_17343# pfet$367
Xpfet$374_3 vdd vdd m1_n4978_24224# vss pfet$374
Xnfet$377_11 m1_27031_17343# vss m1_27190_17836# vss nfet$377
Xpfet$353_8 vdd vdd m1_28113_15778# m1_28470_16080# pfet$353
Xpfet$372_0 vdd vdd m1_n8625_26174# m1_n9336_24346# pfet$372
Xpfet$349_95 vdd vdd m1_21564_17714# m1_22034_17714# pfet$349
Xpfet$349_84 vdd vdd m1_17381_17714# m1_17851_17714# pfet$349
Xpfet$349_73 vdd vdd m1_16538_15778# m1_13668_17714# pfet$349
Xpfet$349_62 vdd vdd m1_23007_17836# m1_22848_17343# pfet$349
Xpfet$349_40 vdd m1_10560_16202# m1_10075_17518# m1_10458_17836# pfet$349
Xpfet$349_51 vdd vdd m1_n1168_15778# m1_n811_16080# pfet$349
Xpfet$351_5 vdd vdd vdd m1_n695_19850# m1_1103_20152# m1_1103_20152# pfet$351
Xnfet$400_0 m1_n7186_25858# vss m1_n7320_25516# vss nfet$400
Xpfet$351_30 vdd vdd vdd m1_24560_19550# m1_21880_15478# m1_21880_15478# pfet$351
Xnfet$374_12 m1_14556_21786# vss m1_15188_21786# vss nfet$374
Xnfet$390_11 m1_15171_20152# m1_15171_20152# m1_n3822_21786# m1_n3822_21786# m1_14005_20470#
+ vss nfet$390
Xnfet$369_23 m1_25424_24346# m1_25424_24346# m1_24309_25858# m1_24309_25858# m1_26371_25502#
+ vss nfet$369
Xnfet$369_12 m1_17058_24346# m1_17058_24346# m1_15943_25858# m1_15943_25858# m1_18005_25502#
+ vss nfet$369
Xnfet$398_0 m1_n9952_24224# m1_n9952_24224# m1_n10308_24542# m1_n10308_24542# m1_n9854_24542#
+ vss nfet$398
Xnfet$371_13 m1_16452_21590# m1_16452_21590# m1_17939_22513# m1_17939_22513# m1_16911_21586#
+ vss nfet$371
Xnfet$377_5 m1_n7247_17714# vss m1_n6657_17518# vss nfet$377
Xnfet$375_2 m1_n7401_15478# vss m1_1103_20152# vss nfet$375
Xnfet$382_3 m1_7522_21786# m1_7522_21786# vss vss m1_6360_21586# vss nfet$382
Xnfet$382_12 m1_18073_21786# m1_18073_21786# vss vss m1_16911_21586# vss nfet$382
Xpfet$367_3 vdd m1_n6172_16202# m1_n6657_17518# m1_n6274_17836# pfet$367
Xpfet$374_4 vdd vdd m1_n5571_25662# m1_n10452_25858# pfet$374
Xnfet$377_12 m1_28470_16080# vss m1_28113_15778# vss nfet$377
Xpfet$353_9 vdd vdd m1_29087_15778# m1_26217_17714# pfet$353
Xnfet$380_0 pd1 vss m1_n1263_21786# vss nfet$380
Xpfet$365_0 vdd m1_32818_20470# m1_32818_20470# m1_33050_19550# m1_30256_19792# m1_30256_19792#
+ pfet$365
Xpfet$372_1 vdd m1_n8625_26174# vdd m1_n8848_25658# pfet$372
Xpfet$349_96 vdd vdd m1_18665_17343# m1_21564_17714# pfet$349
Xpfet$349_85 vdd m1_18926_16202# m1_18441_17518# m1_18824_17836# pfet$349
Xpfet$349_74 vdd vdd m1_14641_17836# m1_14482_17343# pfet$349
Xpfet$349_63 vdd m1_23930_15778# m1_23109_16202# m1_22848_17343# pfet$349
Xpfet$349_30 vdd vdd m1_1933_17343# m1_4832_17714# pfet$349
Xpfet$349_41 vdd vdd m1_10075_17518# m1_9485_17714# pfet$349
Xpfet$349_52 vdd m1_n3064_17714# vdd m1_n1989_16202# pfet$349
Xnfet$400_1 m1_n6856_24542# vss m1_n6111_25858# vss nfet$400
Xpfet$351_6 vdd vdd vdd m1_6339_19850# m1_8137_20152# m1_8137_20152# pfet$351
Xpfet$351_31 vdd m1_n2543_20130# m1_n2543_20130# m1_20407_19850# m1_19969_19550# m1_19969_19550#
+ pfet$351
Xpfet$351_20 vdd m1_n3822_21786# m1_n3822_21786# m1_14009_19550# m1_9015_17714# m1_9015_17714#
+ pfet$351
Xnfet$374_13 m1_16322_21786# vss m1_16452_21590# vss nfet$374
Xnfet$390_12 m1_18688_20152# m1_18688_20152# m1_n1927_20274# m1_n1927_20274# m1_17522_20470#
+ vss nfet$390
Xnfet$369_24 m1_30095_25658# m1_30095_25658# vss vss m1_30554_25502# vss nfet$369
Xnfet$369_13 m1_13363_25658# m1_13363_25658# vss vss m1_13822_25502# vss nfet$369
Xnfet$398_1 m1_n9336_24346# m1_n9336_24346# m1_n8625_26174# m1_n8625_26174# m1_n8389_25502#
+ vss nfet$398
Xnfet$371_14 m1_12805_21786# m1_12805_21786# m1_14422_22513# m1_14422_22513# m1_14026_21586#
+ vss nfet$371
Xnfet$377_6 m1_n7247_17714# vss m1_n7383_17599# vss nfet$377
Xnfet$382_4 m1_1120_21786# m1_1120_21786# vss vss m1_n42_21586# vss nfet$382
Xnfet$382_13 m1_18705_21786# m1_18705_21786# vss vss m1_17543_21586# vss nfet$382
Xpfet$367_4 vdd m1_28113_15778# m1_27292_16202# m1_27031_17343# pfet$367
Xnfet$375_3 m1_649_17714# vss m1_5901_19550# vss nfet$375
Xpfet$374_5 vdd vdd m1_n4847_25662# m1_n10452_25858# pfet$374
Xnfet$377_13 m1_26217_17714# vss m1_25747_17714# vss nfet$377
Xnfet$380_1 pd2 vss m1_2254_21786# vss nfet$380
Xnfet$373_0 m1_9485_17714# vss m1_9015_17714# vss nfet$373
Xpfet$358_0 vdd vdd vdd m1_33050_22344# m1_31535_22102# m1_31535_22102# pfet$358
Xpfet$365_1 vdd vdd vdd m1_33050_19550# m1_31535_19792# m1_31535_19792# pfet$365
Xpfet$372_2 vdd m1_n3651_26174# vdd m1_n4978_24224# pfet$372
Xpfet$349_97 vdd vdd m1_22493_16080# m1_n7513_20152# pfet$349
Xpfet$349_86 vdd m1_19637_18030# vdd m1_18310_16080# pfet$349
Xpfet$349_75 vdd vdd m1_17697_15478# sd3 pfet$349
Xpfet$349_64 vdd vdd m1_23930_15778# m1_24287_16080# pfet$349
Xpfet$349_20 vdd vdd m1_1119_17714# m1_1578_16080# pfet$349
Xpfet$349_31 vdd m1_3372_16080# m1_2905_18030# m1_1933_17343# pfet$349
Xpfet$349_42 vdd m1_11271_18030# vdd m1_9944_16080# pfet$349
Xpfet$349_53 vdd vdd m1_n3218_15478# sd8 pfet$349
Xpfet$351_7 vdd vdd vdd m1_6975_19550# m1_965_15478# m1_965_15478# pfet$351
Xpfet$351_32 vdd m1_n2543_20130# m1_n2543_20130# m1_21043_19550# m1_17381_17714# m1_17381_17714#
+ pfet$351
Xpfet$351_21 vdd vdd vdd m1_13373_19850# m1_15171_20152# m1_15171_20152# pfet$351
Xpfet$351_10 vdd vdd vdd m1_9856_19850# m1_11654_20152# m1_11654_20152# pfet$351
Xnfet$374_14 m1_19839_21786# vss m1_19969_21590# vss nfet$374
Xnfet$390_13 m1_13514_15478# m1_13514_15478# m1_n1927_20274# m1_n1927_20274# m1_16890_20470#
+ vss nfet$390
Xnfet$369_25 m1_29607_24346# m1_29607_24346# m1_28492_25858# m1_28492_25858# m1_30554_25502#
+ vss nfet$369
Xnfet$369_14 m1_12875_24346# m1_12875_24346# m1_11760_25858# m1_11760_25858# m1_13822_25502#
+ vss nfet$369
Xnfet$398_2 m1_n8848_25658# m1_n8848_25658# vss vss m1_n8389_25502# vss nfet$398
Xnfet$377_7 m1_26217_17714# vss m1_26807_17518# vss nfet$377
Xnfet$371_15 m1_26873_21786# m1_26873_21786# m1_28490_22513# m1_28490_22513# m1_28094_21586#
+ vss nfet$371
Xpfet$349_110 vdd vdd m1_10458_17836# m1_10299_17343# pfet$349
Xnfet$382_14 m1_15188_21786# m1_15188_21786# vss vss m1_14026_21586# vss nfet$382
Xpfet$367_5 vdd m1_29087_15778# m1_28470_16080# m1_27190_17836# pfet$367
Xnfet$375_4 m1_4832_17714# vss m1_9418_19550# vss nfet$375
Xpfet$374_6 vdd vdd m1_n4623_25487# fin pfet$374
Xnfet$382_5 m1_4005_21786# m1_4005_21786# vss vss m1_2843_21586# vss nfet$382
Xnfet$380_2 pd9 vss m1_26873_21786# vss nfet$380
Xpfet$354_10 vdd vdd m1_29239_20152# m1_26063_15478# pfet$354
Xnfet$373_1 m1_9015_17714# vss m1_6116_17343# vss nfet$373
Xpfet$365_2 vdd m1_32818_21586# m1_32818_21586# m1_33050_22344# m1_30256_22102# m1_30256_22102#
+ pfet$365
Xpfet$372_3 vdd vdd m1_n3651_26174# m1_n3541_23922# pfet$372
Xpfet$349_98 vdd m1_20104_16080# m1_19637_18030# m1_18665_17343# pfet$349
Xpfet$349_87 vdd vdd m1_18310_16080# m1_n7513_20152# pfet$349
Xpfet$349_76 vdd m1_17851_17714# vdd m1_18926_16202# pfet$349
Xpfet$349_65 vdd m1_24904_15778# m1_24287_16080# m1_23007_17836# pfet$349
Xpfet$349_21 vdd vdd m1_965_15478# sd7 pfet$349
Xpfet$349_10 vdd m1_8172_15778# m1_7555_16080# m1_6275_17836# pfet$349
Xpfet$349_32 vdd vdd m1_2905_18030# m1_3015_15778# pfet$349
Xpfet$349_43 vdd vdd m1_11271_18030# m1_11381_15778# pfet$349
Xpfet$349_54 vdd vdd m1_n1278_18030# m1_n1168_15778# pfet$349
Xpfet$351_8 vdd m1_9624_19404# m1_9624_19404# m1_10492_19550# m1_4832_17714# m1_4832_17714#
+ pfet$351
Xpfet$351_33 vdd m1_n3206_20274# m1_n3206_20274# m1_24560_19550# m1_21564_17714# m1_21564_17714#
+ pfet$351
Xpfet$351_22 vdd vdd vdd m1_14009_19550# m1_9331_15478# m1_9331_15478# pfet$351
Xpfet$351_11 vdd vdd vdd m1_10492_19550# m1_5148_15478# m1_5148_15478# pfet$351
Xpfet$370_0 vdd m1_n10309_25662# m1_n10572_23922# m1_n10796_25662# pfet$370
Xnfet$374_15 m1_28624_21786# vss m1_29256_21786# vss nfet$374
Xnfet$390_14 m1_22205_20152# m1_22205_20152# m1_n2543_20130# m1_n2543_20130# m1_21039_20470#
+ vss nfet$390
Xnfet$398_3 m1_n9336_24346# m1_n9336_24346# vss vss m1_n9854_24542# vss nfet$398
Xnfet$369_26 m1_25912_25658# m1_25912_25658# vss vss m1_26371_25502# vss nfet$369
Xnfet$369_15 m1_25424_24346# m1_25424_24346# vss vss m1_24906_24542# vss nfet$369
Xnfet$377_8 m1_n7513_20152# vss m1_26676_16080# vss nfet$377
Xnfet$371_16 m1_27003_21590# m1_27003_21590# m1_28490_22513# m1_28490_22513# m1_27462_21586#
+ vss nfet$371
Xnfet$396_0 m1_n3822_20130# m1_n3822_20130# m1_n4485_20152# m1_n4485_20152# m1_n3724_20470#
+ vss nfet$396
Xpfet$349_100 vdd vdd m1_23820_18030# m1_23930_15778# pfet$349
Xnfet$382_15 m1_14556_21786# m1_14556_21786# vss vss m1_13394_21586# vss nfet$382
Xnfet$375_5 m1_965_15478# vss m1_8137_20152# vss nfet$375
Xnfet$382_6 m1_4637_21786# m1_4637_21786# vss vss m1_3475_21586# vss nfet$382
Xpfet$367_6 vdd m1_28470_16080# m1_28003_18030# m1_27031_17343# pfet$367
Xpfet$374_7 vdd vdd m1_n3541_23922# m1_n3184_24224# pfet$374
Xpfet$354_11 vdd vdd m1_18688_20152# m1_13514_15478# pfet$354
Xnfet$373_2 m1_6275_17836# m1_7555_16080# m1_7088_18030# vss nfet$373
Xpfet$372_4 vdd m1_n10452_25858# vdd m1_n4362_24346# pfet$372
Xpfet$349_99 vdd m1_23109_16202# m1_22624_17518# m1_23007_17836# pfet$349
Xpfet$349_88 vdd vdd m1_18441_17518# m1_17851_17714# pfet$349
Xpfet$349_77 vdd vdd m1_17851_17714# m1_18310_16080# pfet$349
Xpfet$349_66 vdd vdd m1_24904_15778# m1_22034_17714# pfet$349
Xpfet$349_22 vdd vdd m1_3015_15778# m1_3372_16080# pfet$349
Xpfet$349_11 vdd vdd m1_9485_17714# m1_9944_16080# pfet$349
Xpfet$349_33 vdd vdd m1_5892_17518# m1_5302_17714# pfet$349
Xpfet$349_44 vdd vdd m1_649_17714# m1_1119_17714# pfet$349
Xpfet$349_55 vdd vdd m1_n2474_17518# m1_n3064_17714# pfet$349
Xpfet$351_9 vdd m1_9624_19404# m1_9624_19404# m1_9856_19850# m1_9418_19550# m1_9418_19550#
+ pfet$351
Xpfet$363_0 vdd vdd vdd m1_36073_22344# define define pfet$363
Xpfet$351_34 vdd m1_n3206_20274# m1_n3206_20274# m1_23924_19850# m1_23486_19550# m1_23486_19550#
+ pfet$351
Xpfet$351_23 vdd vdd vdd m1_16890_19850# m1_18688_20152# m1_18688_20152# pfet$351
Xpfet$351_12 vdd m1_6107_19404# m1_6107_19404# m1_6975_19550# m1_649_17714# m1_649_17714#
+ pfet$351
Xpfet$370_1 vdd m1_n9952_24224# m1_n8848_25658# m1_n10933_25858# pfet$370
Xnfet$374_16 m1_26873_21786# vss m1_27003_21590# vss nfet$374
Xnfet$390_15 m1_17697_15478# m1_17697_15478# m1_n2543_20130# m1_n2543_20130# m1_20407_20470#
+ vss nfet$390
Xnfet$369_27 m1_12875_24346# m1_12875_24346# vss vss m1_12357_24542# vss nfet$369
Xnfet$369_16 m1_24808_24224# m1_24808_24224# m1_24452_24542# m1_24452_24542# m1_24906_24542#
+ vss nfet$369
Xnfet$398_4 m1_n4978_24224# m1_n4978_24224# m1_n10452_25858# m1_n10452_25858# m1_n4880_24542#
+ vss nfet$398
Xnfet$377_9 m1_n10452_25858# vss m1_27031_17343# vss nfet$377
Xnfet$371_17 m1_12935_21590# m1_12935_21590# m1_14422_22513# m1_14422_22513# m1_13394_21586#
+ vss nfet$371
Xnfet$389_0 m1_7198_15778# m1_7198_15778# m1_7088_18030# m1_7088_18030# m1_7324_17358#
+ vss nfet$389
Xnfet$396_1 m1_n1927_20274# m1_n1927_20274# vss vss m1_n2445_20470# vss nfet$396
Xpfet$349_101 vdd vdd m1_19637_18030# m1_19747_15778# pfet$349
Xnfet$382_7 m1_488_21786# m1_488_21786# vss vss m1_n674_21586# vss nfet$382
Xnfet$375_6 m1_9015_17714# vss m1_12935_19550# vss nfet$375
Xnfet$382_16 m1_28624_21786# m1_28624_21786# vss vss m1_27462_21586# vss nfet$382
Xpfet$367_7 vdd m1_27292_16202# m1_26807_17518# m1_27190_17836# pfet$367
Xpfet$374_8 vdd vdd m1_n2567_23922# m1_n7320_25516# pfet$374
Xpfet$354_12 vdd vdd m1_15171_20152# m1_9331_15478# pfet$354
Xnfet$373_3 m1_n7513_20152# vss m1_9944_16080# vss nfet$373
Xpfet$372_5 vdd vdd m1_n10308_24542# m1_n9952_24224# pfet$372
Xpfet$349_89 vdd vdd m1_22848_17343# m1_25747_17714# pfet$349
Xpfet$349_78 vdd vdd m1_13514_15478# sd4 pfet$349
Xpfet$349_67 vdd m1_22034_17714# vdd m1_23109_16202# pfet$349
Xpfet$349_12 vdd m1_3989_15778# m1_3372_16080# m1_2092_17836# pfet$349
Xpfet$349_23 vdd m1_5302_17714# vdd m1_6377_16202# pfet$349
Xpfet$349_34 vdd vdd m1_5761_16080# m1_n7513_20152# pfet$349
Xpfet$349_45 vdd vdd m1_9944_16080# m1_n7513_20152# pfet$349
Xpfet$349_56 vdd m1_n1278_18030# vdd m1_n2605_16080# pfet$349
Xnfet$371_0 m1_n1133_21590# m1_n1133_21590# m1_354_22513# m1_354_22513# m1_n674_21586#
+ vss nfet$371
Xpfet$363_1 vdd m1_35837_22102# m1_35837_22102# m1_36073_22344# fout fout pfet$363
Xpfet$370_2 vdd m1_n4362_24346# m1_n4847_25662# m1_n4464_25980# pfet$370
Xpfet$356_0 vdd vdd m1_n647_25662# m1_n789_25858# pfet$356
Xpfet$351_35 vdd m1_n3822_21786# m1_n3822_21786# m1_13373_19850# m1_12935_19550# m1_12935_19550#
+ pfet$351
Xpfet$351_24 vdd m1_n1927_20274# m1_n1927_20274# m1_16890_19850# m1_16452_19550# m1_16452_19550#
+ pfet$351
Xpfet$351_13 vdd m1_n927_19404# m1_n927_19404# m1_n695_19850# m1_n1133_19550# m1_n1133_19550#
+ pfet$351
Xnfet$374_17 m1_25107_21786# vss m1_25739_21786# vss nfet$374
Xnfet$390_16 m1_25722_20152# m1_25722_20152# m1_n3206_20274# m1_n3206_20274# m1_24556_20470#
+ vss nfet$390
Xnfet$369_17 m1_20625_24224# m1_20625_24224# m1_20269_24542# m1_20269_24542# m1_20723_24542#
+ vss nfet$369
Xnfet$398_5 m1_n4362_24346# m1_n4362_24346# vss vss m1_n4880_24542# vss nfet$398
Xnfet$389_1 m1_5761_16080# m1_5761_16080# vss vss m1_7324_17358# vss nfet$389
Xnfet$396_2 m1_n3206_20274# m1_n3206_20274# vss vss m1_n3724_20470# vss nfet$396
Xnfet$382_8 m1_25739_21786# m1_25739_21786# vss vss m1_24577_21586# vss nfet$382
Xpfet$349_102 vdd vdd m1_13198_17714# m1_13668_17714# pfet$349
Xnfet$375_7 m1_5148_15478# vss m1_11654_20152# vss nfet$375
Xnfet$382_17 m1_29256_21786# m1_29256_21786# vss vss m1_28094_21586# vss nfet$382
Xpfet$374_9 vdd vdd m1_n4464_25980# m1_n4623_25487# pfet$374
Xpfet$354_13 vdd vdd m1_16452_19550# m1_13198_17714# pfet$354
Xnfet$373_4 m1_10299_17343# m1_10560_16202# m1_10075_17518# vss nfet$373
Xpfet$349_13 vdd vdd m1_5148_15478# sd6 pfet$349
Xpfet$372_6 vdd m1_n10308_24542# vdd m1_n9336_24346# pfet$372
Xpfet$349_79 vdd m1_15564_15778# m1_14743_16202# m1_14482_17343# pfet$349
Xpfet$349_68 vdd vdd m1_22034_17714# m1_22493_16080# pfet$349
Xpfet$349_24 vdd m1_6377_16202# m1_5892_17518# m1_6275_17836# pfet$349
Xpfet$349_35 vdd vdd m1_9015_17714# m1_9485_17714# pfet$349
Xpfet$349_46 vdd vdd m1_n2250_17343# m1_649_17714# pfet$349
Xpfet$349_57 vdd m1_n1989_16202# m1_n2474_17518# m1_n2091_17836# pfet$349
Xpfet$349_0 vdd vdd m1_12355_15778# m1_9485_17714# pfet$349
Xnfet$371_1 m1_n1263_21786# m1_n1263_21786# m1_354_22513# m1_354_22513# m1_n42_21586#
+ vss nfet$371
Xpfet$356_1 vdd vdd m1_n1134_25662# m1_n1271_25858# pfet$356
Xpfet$370_3 vdd m1_n3184_24224# m1_n3651_26174# m1_n4623_25487# pfet$370
Xpfet$351_25 vdd vdd vdd m1_17526_19550# m1_13514_15478# m1_13514_15478# pfet$351
Xpfet$351_14 vdd m1_n927_19404# m1_n927_19404# m1_n59_19550# m1_n7383_17599# m1_n7383_17599#
+ pfet$351
Xnfet$390_17 m1_21880_15478# m1_21880_15478# m1_n3206_20274# m1_n3206_20274# m1_23924_20470#
+ vss nfet$390
Xnfet$369_18 m1_21241_24346# m1_21241_24346# vss vss m1_20723_24542# vss nfet$369
Xnfet$398_6 m1_n4978_24224# m1_n4978_24224# vss vss m1_n3415_25502# vss nfet$398
Xnfet$389_2 m1_9944_16080# m1_9944_16080# vss vss m1_11507_17358# vss nfet$389
Xnfet$396_3 m1_n6973_21481# m1_n6973_21481# m1_n6839_20152# m1_n6839_20152# m1_n6282_20470#
+ vss nfet$396
Xnfet$382_9 m1_25107_21786# m1_25107_21786# vss vss m1_23945_21586# vss nfet$382
Xpfet$349_103 vdd m1_14743_16202# m1_14258_17518# m1_14641_17836# pfet$349
Xnfet$375_8 m1_n7383_17599# vss m1_n1133_19550# vss nfet$375
Xnfet$394_0 m1_n10452_25858# m1_n10452_25858# m1_n7186_25858# m1_n7186_25858# m1_n6629_25502#
+ vss nfet$394
Xpfet$354_14 vdd vdd m1_23486_19550# m1_21564_17714# pfet$354
Xpfet$379_0 vdd vdd vdd m1_n5019_19550# m1_n4485_20152# m1_n4485_20152# pfet$379
Xnfet$373_5 m1_10458_17836# m1_11738_16080# m1_11271_18030# vss nfet$373
Xpfet$372_7 vdd vdd m1_n10452_25858# m1_n4978_24224# pfet$372
Xpfet$349_69 vdd vdd m1_20721_15778# m1_17851_17714# pfet$349
Xpfet$349_14 vdd vdd m1_2092_17836# m1_1933_17343# pfet$349
Xpfet$349_25 vdd vdd m1_1709_17518# m1_1119_17714# pfet$349
Xpfet$349_36 vdd vdd m1_6116_17343# m1_9015_17714# pfet$349
Xpfet$349_47 vdd m1_11738_16080# m1_11271_18030# m1_10299_17343# pfet$349
Xpfet$349_58 vdd vdd m1_n3534_17714# m1_n3064_17714# pfet$349
Xpfet$370_4 vdd m1_n2567_23922# m1_n3184_24224# m1_n4464_25980# pfet$370
Xnfet$371_2 m1_9288_21786# m1_9288_21786# m1_9645_21447# m1_9645_21447# m1_10509_21586#
+ vss nfet$371
Xpfet$351_26 vdd m1_n1927_20274# m1_n1927_20274# m1_17526_19550# m1_13198_17714# m1_13198_17714#
+ pfet$351
Xpfet$351_15 vdd vdd vdd m1_n59_19550# m1_n7401_15478# m1_n7401_15478# pfet$351
Xpfet$349_1 vdd vdd m1_11381_15778# m1_11738_16080# pfet$349
Xpfet$356_2 vdd vdd m1_n1271_25858# m1_n10452_25858# pfet$356
Xpfet$361_0 vdd vdd m1_n1263_21786# pd1 pfet$361
Xnfet$369_19 m1_21729_25658# m1_21729_25658# vss vss m1_22188_25502# vss nfet$369
Xnfet$398_7 m1_n3541_23922# m1_n3541_23922# m1_n3651_26174# m1_n3651_26174# m1_n3415_25502#
+ vss nfet$398
Xnfet$389_3 m1_11381_15778# m1_11381_15778# m1_11271_18030# m1_11271_18030# m1_11507_17358#
+ vss nfet$389
Xnfet$396_4 m1_2590_19404# m1_2590_19404# vss vss m1_n2445_21430# vss nfet$396
Xpfet$349_104 vdd vdd m1_14127_16080# m1_n7513_20152# pfet$349
Xnfet$375_9 m1_25747_17714# vss m1_27003_19550# vss nfet$375
Xnfet$394_1 m1_n6111_25858# m1_n6111_25858# vss vss m1_n6629_25502# vss nfet$394
Xnfet$387_0 m1_34093_22102# vss fout vss nfet$387
Xpfet$354_15 vdd vdd m1_22205_20152# m1_17697_15478# pfet$354
Xnfet$373_6 m1_6116_17343# vss m1_6275_17836# vss nfet$373
Xpfet$349_15 vdd vdd m1_5302_17714# m1_5761_16080# pfet$349
Xpfet$349_26 vdd vdd m1_4832_17714# m1_5302_17714# pfet$349
Xpfet$349_37 vdd m1_7555_16080# m1_7088_18030# m1_6116_17343# pfet$349
Xpfet$349_48 vdd vdd m1_n3064_17714# m1_n2605_16080# pfet$349
Xpfet$349_59 vdd vdd m1_n2605_16080# m1_n7513_20152# pfet$349
Xnfet$371_3 m1_9418_21590# m1_9418_21590# m1_9645_21447# m1_9645_21447# m1_9877_21586#
+ vss nfet$371
Xpfet$351_27 vdd vdd vdd m1_20407_19850# m1_22205_20152# m1_22205_20152# pfet$351
Xpfet$351_16 vdd vdd vdd m1_28077_19550# m1_26063_15478# m1_26063_15478# pfet$351
Xpfet$356_3 vdd vdd m1_1607_24542# m1_n789_25858# pfet$356
Xpfet$349_2 vdd m1_12355_15778# m1_11738_16080# m1_10458_17836# pfet$349
Xpfet$370_5 vdd m1_n10572_23922# m1_n10308_24542# m1_n10933_25858# pfet$370
Xpfet$361_1 vdd vdd m1_2254_21786# pd2 pfet$361
Xpfet$354_0 vdd vdd m1_2384_19550# m1_n3534_17714# pfet$354
Xnfet$389_4 m1_10560_16202# m1_10560_16202# vss vss m1_10042_16398# vss nfet$389
Xnfet$396_5 m1_6107_19404# m1_6107_19404# m1_n5227_21418# m1_n5227_21418# m1_n2445_21430#
+ vss nfet$396
Xpfet$349_105 vdd vdd m1_14258_17518# m1_13668_17714# pfet$349
Xpfet$354_16 vdd vdd m1_19969_19550# m1_17381_17714# pfet$354
Xnfet$373_7 m1_9485_17714# vss m1_10075_17518# vss nfet$373
Xpfet$349_16 vdd vdd m1_3989_15778# m1_1119_17714# pfet$349
Xpfet$349_27 vdd m1_2194_16202# m1_1709_17518# m1_2092_17836# pfet$349
Xpfet$349_38 vdd vdd m1_7088_18030# m1_7198_15778# pfet$349
Xpfet$349_49 vdd m1_n194_15778# m1_n811_16080# m1_n2091_17836# pfet$349
Xnfet$371_4 m1_5901_21590# m1_5901_21590# m1_7388_22513# m1_7388_22513# m1_6360_21586#
+ vss nfet$371
Xpfet$351_28 vdd vdd vdd m1_21043_19550# m1_17697_15478# m1_17697_15478# pfet$351
Xpfet$351_17 vdd m1_n3822_20130# m1_n3822_20130# m1_28077_19550# m1_25747_17714# m1_25747_17714#
+ pfet$351
Xpfet$356_4 vdd vdd m1_488_21786# m1_n789_25858# pfet$356
Xpfet$349_3 vdd m1_11381_15778# m1_10560_16202# m1_10299_17343# pfet$349
Xpfet$370_6 vdd m1_n8848_25658# m1_n8055_24542# m1_n10796_25662# pfet$370
Xpfet$361_2 vdd vdd m1_26873_21786# pd9 pfet$361
Xpfet$354_1 vdd vdd m1_4620_20152# m1_n3218_15478# pfet$354
Xnfet$389_5 m1_9944_16080# m1_9944_16080# m1_9485_17714# m1_9485_17714# m1_10042_16398#
+ vss nfet$389
Xnfet$396_6 m1_n5764_21786# m1_n5764_21786# vss vss m1_n6282_21430# vss nfet$396
Xpfet$349_106 vdd vdd m1_14482_17343# m1_17381_17714# pfet$349
Xpfet$354_17 vdd vdd m1_25722_20152# m1_21880_15478# pfet$354
Xnfet$372_10 m1_9015_17714# m1_9015_17714# vss vss m1_14005_20470# vss nfet$372
Xnfet$373_8 m1_7555_16080# vss m1_7198_15778# vss nfet$373
Xnfet$392_0 m1_n6274_17836# m1_n4994_16080# m1_n5461_18030# vss nfet$392
Xpfet$349_17 vdd vdd m1_n2091_17836# m1_n2250_17343# pfet$349
Xpfet$349_28 vdd m1_2905_18030# vdd m1_1578_16080# pfet$349
Xpfet$349_39 vdd m1_7088_18030# vdd m1_5761_16080# pfet$349
Xpfet$377_0 vdd m1_n6380_21786# m1_n6380_21786# m1_n5019_19550# m1_n5227_20152# m1_n5227_20152#
+ pfet$377
Xnfet$371_5 m1_2254_21786# m1_2254_21786# m1_3871_22513# m1_3871_22513# m1_3475_21586#
+ vss nfet$371
Xpfet$356_5 vdd vdd m1_326_24346# m1_n7513_20152# pfet$356
Xpfet$349_4 vdd m1_9485_17714# vdd m1_10560_16202# pfet$349
Xnfet$405_0 m1_n6839_20152# vss m1_n8145_21908# vss nfet$405
Xpfet$370_7 vdd m1_n3541_23922# m1_n4362_24346# m1_n4623_25487# pfet$370
Xpfet$351_29 vdd vdd vdd m1_23924_19850# m1_25722_20152# m1_25722_20152# pfet$351
Xpfet$351_18 vdd vdd vdd m1_27441_19850# m1_29239_20152# m1_29239_20152# pfet$351
Xpfet$354_2 vdd vdd m1_1103_20152# m1_n7401_15478# pfet$354
Xnfet$375_10 m1_26063_15478# vss m1_29239_20152# vss nfet$375
Xnfet$389_6 m1_1578_16080# m1_1578_16080# vss vss m1_3141_17358# vss nfet$389
Xnfet$396_7 m1_n3822_21786# m1_n3822_21786# m1_n4485_21904# m1_n4485_21904# m1_n3724_21430#
+ vss nfet$396
Xpfet$349_107 vdd m1_15921_16080# m1_15454_18030# m1_14482_17343# pfet$349
Xnfet$372_11 m1_13198_17714# m1_13198_17714# vss vss m1_17522_20470# vss nfet$372
Xnfet$373_9 sd5 vss m1_9331_15478# vss nfet$373
Xnfet$385_0 m1_31535_22102# m1_32818_21586# vss vss nfet$385
Xpfet$349_18 vdd m1_1119_17714# vdd m1_2194_16202# pfet$349
Xnfet$392_1 m1_n6433_17343# m1_n4377_15778# m1_n4994_16080# vss nfet$392
Xpfet$377_1 vdd vdd vdd m1_n5019_22344# m1_n4485_21904# m1_n4485_21904# pfet$377
Xpfet$349_29 vdd vdd m1_1578_16080# m1_n7513_20152# pfet$349
.ends

.subckt nfet$440 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$416 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$414 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$441 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$417 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$415 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$439 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$442 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_drive_buffer$5 vss in vdd out
Xnfet$440_0 out out vss m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# m1_4274_n1060#
+ m1_4274_n1060# out m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# vss vss
+ nfet$440
Xpfet$416_0 vdd vdd m1_4002_n1060# m1_3466_n454# pfet$416
Xpfet$414_0 out out m1_4274_n1060# vdd m1_4274_n1060# out vdd vdd m1_4274_n1060# out
+ m1_4274_n1060# m1_4274_n1060# out m1_4274_n1060# vdd m1_4274_n1060# vdd m1_4274_n1060#
+ pfet$414
Xnfet$441_0 m1_3466_n454# vss m1_4002_n1060# vss nfet$441
Xpfet$417_0 vdd vdd m1_3466_n454# in pfet$417
Xpfet$415_0 m1_4274_n1060# vdd vdd m1_4274_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ vdd m1_4002_n1060# m1_4002_n1060# pfet$415
Xnfet$439_0 m1_4274_n1060# vss m1_4002_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ m1_4274_n1060# vss m1_4002_n1060# vss nfet$439
Xnfet$442_0 in vss m1_3466_n454# vss nfet$442
.ends

.subckt nfet$410 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$385 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt inv1u05u$3 VDD in VSS out
Xnfet$410_0 in VSS out VSS nfet$410
Xpfet$385_0 VDD VDD out in pfet$385
.ends

.subckt pfet$381 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_954_0# w_n180_n88# a_854_n136#
+ a_n92_0# a_446_n136# a_650_n136# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt nfet$409 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$384 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pass1u05u$3 VDD VSS ind ins clkn clkp
Xnfet$409_0 clkn ind ins VSS nfet$409
Xpfet$384_0 VDD ind ins clkp pfet$384
.ends

.subckt nfet$407 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$382 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_954_0# w_n180_n88#
+ a_38_n60# a_n92_0# a_1058_n60# a_854_n60# a_342_0# a_138_0# a_650_n60#
X0 a_954_0# a_854_n60# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n60# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt nfet$406 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt nfet$408 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$383 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=4.55p ps=15.3u w=7u l=0.5u
.ends

.subckt nfet$411 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$386 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.5u
.ends

.subckt xp_programmable_basic_pump$2 up vdd s1 s2 s3 s4 down out iref vss
Xinv1u05u$3_2 vdd s2 vss inv1u05u$3_2/out inv1u05u$3
Xpfet$381_17 m1_n8156_628# m1_n8156_628# pass1u05u$3_7/ins out out vdd pass1u05u$3_7/ins
+ m1_n8156_628# pass1u05u$3_7/ins pass1u05u$3_7/ins m1_n8156_628# out pass1u05u$3_7/ins
+ pass1u05u$3_7/ins pfet$381
Xpass1u05u$3_6 vdd vss iref pass1u05u$3_6/ins s4 inv1u05u$3_0/out pass1u05u$3
Xnfet$407_5 vss vss vss vss vss vss nfet$407
Xpfet$382_0 vdd vdd m1_n4127_3649# vss vss m1_n4127_3649# vdd vss vdd vss vss vdd
+ m1_n4127_3649# vss pfet$382
Xinv1u05u$3_3 vdd s1 vss inv1u05u$3_3/out inv1u05u$3
Xpfet$381_18 m1_n8156_628# m1_n8156_628# pass1u05u$3_7/ins out out vdd pass1u05u$3_7/ins
+ m1_n8156_628# pass1u05u$3_7/ins pass1u05u$3_7/ins m1_n8156_628# out pass1u05u$3_7/ins
+ pass1u05u$3_7/ins pfet$381
Xpass1u05u$3_7 vdd vss pass1u05u$3_7/ind pass1u05u$3_7/ins s4 inv1u05u$3_0/out pass1u05u$3
Xnfet$407_6 down down vss vss m1_n8807_n11192# vss nfet$407
Xpfet$382_1 m1_n5580_883# m1_n5580_883# out pass1u05u$3_5/ins pass1u05u$3_5/ins out
+ vdd pass1u05u$3_5/ins m1_n5580_883# pass1u05u$3_5/ins pass1u05u$3_5/ins m1_n5580_883#
+ out pass1u05u$3_5/ins pfet$382
Xpfet$381_19 m1_n8156_628# m1_n8156_628# pass1u05u$3_7/ins out out vdd pass1u05u$3_7/ins
+ m1_n8156_628# pass1u05u$3_7/ins pass1u05u$3_7/ins m1_n8156_628# out pass1u05u$3_7/ins
+ pass1u05u$3_7/ins pfet$381
Xnfet$407_7 down down vss vss m1_n8807_n11192# vss nfet$407
Xpfet$382_2 m1_n5580_883# m1_n5580_883# out pass1u05u$3_5/ins pass1u05u$3_5/ins out
+ vdd pass1u05u$3_5/ins m1_n5580_883# pass1u05u$3_5/ins pass1u05u$3_5/ins m1_n5580_883#
+ out pass1u05u$3_5/ins pfet$382
Xnfet$407_8 down down vss vss m1_n8807_n11192# vss nfet$407
Xpfet$382_3 m1_n5580_883# m1_n5580_883# out pass1u05u$3_5/ins pass1u05u$3_5/ins out
+ vdd pass1u05u$3_5/ins m1_n5580_883# pass1u05u$3_5/ins pass1u05u$3_5/ins m1_n5580_883#
+ out pass1u05u$3_5/ins pfet$382
Xnfet$407_9 down down vss vss m1_n8807_n11192# vss nfet$407
Xpfet$382_4 m1_n5580_883# m1_n5580_883# out pass1u05u$3_5/ins pass1u05u$3_5/ins out
+ vdd pass1u05u$3_5/ins m1_n5580_883# pass1u05u$3_5/ins pass1u05u$3_5/ins m1_n5580_883#
+ out pass1u05u$3_5/ins pfet$382
Xnfet$406_10 pass1u05u$3_2/ins pass1u05u$3_2/ins m1_n7679_n8960# m1_n7679_n8960# out
+ vss nfet$406
Xpfet$382_5 m1_n4127_3649# m1_n4127_3649# pass1u05u$3_7/ind pass1u05u$3_7/ind pass1u05u$3_7/ind
+ pass1u05u$3_7/ind vdd pass1u05u$3_7/ind m1_n4127_3649# pass1u05u$3_7/ind pass1u05u$3_7/ind
+ m1_n4127_3649# pass1u05u$3_7/ind pass1u05u$3_7/ind pfet$382
Xnfet$406_11 vss vss vss vss vss vss nfet$406
Xnfet$406_12 down down vss vss m1_n7679_n8960# vss nfet$406
Xnfet$406_13 vss vss vss vss vss vss nfet$406
Xnfet$406_14 vss vss vss vss vss vss nfet$406
Xnfet$406_15 vss vss vss vss vss vss nfet$406
Xnfet$408_0 m1_n7879_n12170# pass1u05u$3_0/ins m1_n7879_n12170# out pass1u05u$3_0/ins
+ vss nfet$408
Xnfet$408_1 m1_n7879_n12170# pass1u05u$3_0/ins m1_n7879_n12170# out pass1u05u$3_0/ins
+ vss nfet$408
Xnfet$408_2 vss down vss m1_n7879_n12170# down vss nfet$408
Xnfet$406_0 pass1u05u$3_6/ins pass1u05u$3_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$406
Xnfet$408_3 vss down vss m1_n7879_n12170# down vss nfet$408
Xnfet$408_4 vss down vss m1_n7879_n12170# down vss nfet$408
Xnfet$406_1 pass1u05u$3_6/ins pass1u05u$3_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$406
Xpfet$383_20 vdd vdd vdd vdd pfet$383
Xnfet$408_5 vss down vss m1_n7879_n12170# down vss nfet$408
Xnfet$411_0 inv1u05u$3_2/out pass1u05u$3_1/ins vss vss nfet$411
Xnfet$406_2 pass1u05u$3_6/ins pass1u05u$3_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$406
Xpfet$383_0 vdd vdd vdd vdd pfet$383
Xnfet$407_10 vss vss vss vss vss vss nfet$407
Xnfet$408_6 m1_n7879_n12170# pass1u05u$3_0/ins m1_n7879_n12170# out pass1u05u$3_0/ins
+ vss nfet$408
Xpfet$383_21 vdd vdd vdd vdd pfet$383
Xnfet$406_3 vss vss vss vss vss vss nfet$406
Xpfet$383_1 vdd vdd vdd vdd pfet$383
Xpfet$383_10 vdd vdd vdd vdd pfet$383
Xnfet$411_1 inv1u05u$3_3/out pass1u05u$3_2/ins vss vss nfet$411
Xnfet$407_11 vss vss vss vss vss vss nfet$407
Xnfet$408_7 m1_n7879_n12170# pass1u05u$3_0/ins m1_n7879_n12170# out pass1u05u$3_0/ins
+ vss nfet$408
Xpfet$383_22 vdd vdd vdd vdd pfet$383
Xnfet$411_2 inv1u05u$3_0/out pass1u05u$3_6/ins vss vss nfet$411
Xnfet$406_4 pass1u05u$3_6/ins pass1u05u$3_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$406
Xpfet$383_2 vdd vdd vdd vdd pfet$383
Xpfet$383_11 vdd vdd vdd vdd pfet$383
Xnfet$407_12 vss vss vss vss vss vss nfet$407
Xpfet$383_23 vdd vdd vdd vdd pfet$383
Xnfet$406_5 vss vss vss vss vss vss nfet$406
Xnfet$408_8 vss vdd vss m1_n8144_n9165# vdd vss nfet$408
Xpfet$383_3 vdd vdd vdd vdd pfet$383
Xpfet$383_12 vdd vdd vdd vdd pfet$383
Xnfet$411_3 inv1u05u$3_1/out pass1u05u$3_0/ins vss vss nfet$411
Xpfet$381_0 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$381
Xnfet$407_13 vss vss vss vss vss vss nfet$407
Xnfet$408_9 m1_n7216_n8262# iref m1_n7216_n8262# pass1u05u$3_7/ind iref vss nfet$408
Xpfet$383_13 vdd vdd vdd vdd pfet$383
Xnfet$406_6 pass1u05u$3_6/ins pass1u05u$3_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$406
Xpfet$383_4 vdd vdd vdd vdd pfet$383
Xpfet$381_1 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$381
Xpfet$383_14 vdd vdd vdd vdd pfet$383
Xnfet$406_7 pass1u05u$3_6/ins pass1u05u$3_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$406
Xpfet$381_2 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$381
Xpfet$383_5 vdd vdd vdd vdd pfet$383
Xpfet$383_15 vdd vdd vdd vdd pfet$383
Xnfet$406_8 pass1u05u$3_6/ins pass1u05u$3_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$406
Xpfet$383_6 vdd vdd vdd vdd pfet$383
Xpfet$381_3 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$381
Xpfet$383_16 vdd vdd vdd vdd pfet$383
Xnfet$406_9 pass1u05u$3_6/ins pass1u05u$3_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$406
Xpfet$381_4 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$381
Xpfet$383_7 vdd vdd vdd vdd pfet$383
Xpfet$383_17 vdd vdd vdd vdd pfet$383
Xpfet$383_8 vdd vdd vdd vdd pfet$383
Xpfet$381_5 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$381
Xpfet$383_18 vdd vdd vdd vdd pfet$383
Xpfet$381_6 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$381
Xpfet$383_9 vdd vdd vdd vdd pfet$383
Xpfet$383_19 vdd vdd vdd vdd pfet$383
Xpfet$381_7 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$381
Xpfet$381_8 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$381
Xpfet$381_20 m1_n8156_628# m1_n8156_628# pass1u05u$3_7/ins out out vdd pass1u05u$3_7/ins
+ m1_n8156_628# pass1u05u$3_7/ins pass1u05u$3_7/ins m1_n8156_628# out pass1u05u$3_7/ins
+ pass1u05u$3_7/ins pfet$381
Xpfet$381_9 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$381
Xpfet$381_21 m1_n6703_2564# m1_n6703_2564# pass1u05u$3_4/ins out out vdd pass1u05u$3_4/ins
+ m1_n6703_2564# pass1u05u$3_4/ins pass1u05u$3_4/ins m1_n6703_2564# out pass1u05u$3_4/ins
+ pass1u05u$3_4/ins pfet$381
Xpfet$381_10 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$381
Xnfet$408_10 m1_n8607_n8040# pass1u05u$3_1/ins m1_n8607_n8040# out pass1u05u$3_1/ins
+ vss nfet$408
Xpass1u05u$3_0 vdd vss iref pass1u05u$3_0/ins s3 inv1u05u$3_1/out pass1u05u$3
Xpfet$386_0 vdd s3 pass1u05u$3_5/ins vdd pfet$386
Xpfet$381_22 m1_n8156_628# m1_n8156_628# pass1u05u$3_7/ins out out vdd pass1u05u$3_7/ins
+ m1_n8156_628# pass1u05u$3_7/ins pass1u05u$3_7/ins m1_n8156_628# out pass1u05u$3_7/ins
+ pass1u05u$3_7/ins pfet$381
Xpfet$381_11 vdd vdd up m1_n5450_4559# m1_n5450_4559# vdd up vdd up up vdd m1_n5450_4559#
+ up up pfet$381
Xnfet$408_11 m1_n8144_n9165# iref m1_n8144_n9165# iref iref vss nfet$408
Xpfet$386_1 vdd s2 pass1u05u$3_4/ins vdd pfet$386
Xpfet$381_23 m1_n8156_628# m1_n8156_628# pass1u05u$3_7/ins out out vdd pass1u05u$3_7/ins
+ m1_n8156_628# pass1u05u$3_7/ins pass1u05u$3_7/ins m1_n8156_628# out pass1u05u$3_7/ins
+ pass1u05u$3_7/ins pfet$381
Xpass1u05u$3_1 vdd vss iref pass1u05u$3_1/ins s2 inv1u05u$3_2/out pass1u05u$3
Xnfet$407_0 down down vss vss m1_n8807_n11192# vss nfet$407
Xpfet$381_12 vdd vdd up m1_n6703_2564# m1_n6703_2564# vdd up vdd up up vdd m1_n6703_2564#
+ up up pfet$381
Xnfet$408_12 vss down vss m1_n8607_n8040# down vss nfet$408
Xpass1u05u$3_2 vdd vss iref pass1u05u$3_2/ins s1 inv1u05u$3_3/out pass1u05u$3
Xpfet$386_2 vdd s1 pass1u05u$3_3/ins vdd pfet$386
Xnfet$407_1 down down vss vss m1_n8807_n11192# vss nfet$407
Xpfet$381_24 m1_n5450_4559# m1_n5450_4559# pass1u05u$3_3/ins out out vdd pass1u05u$3_3/ins
+ m1_n5450_4559# pass1u05u$3_3/ins pass1u05u$3_3/ins m1_n5450_4559# out pass1u05u$3_3/ins
+ pass1u05u$3_3/ins pfet$381
Xpfet$381_13 vdd vdd up m1_n6703_2564# m1_n6703_2564# vdd up vdd up up vdd m1_n6703_2564#
+ up up pfet$381
Xnfet$408_13 vss vdd vss m1_n7216_n8262# vdd vss nfet$408
Xpfet$386_3 vdd s4 pass1u05u$3_7/ins vdd pfet$386
Xpfet$381_25 m1_n6703_2564# m1_n6703_2564# pass1u05u$3_4/ins out out vdd pass1u05u$3_4/ins
+ m1_n6703_2564# pass1u05u$3_4/ins pass1u05u$3_4/ins m1_n6703_2564# out pass1u05u$3_4/ins
+ pass1u05u$3_4/ins pfet$381
Xpass1u05u$3_3 vdd vss pass1u05u$3_7/ind pass1u05u$3_3/ins s1 inv1u05u$3_3/out pass1u05u$3
Xnfet$407_2 down down vss vss m1_n8807_n11192# vss nfet$407
Xpfet$381_14 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$381
Xnfet$408_14 m1_n8607_n8040# pass1u05u$3_1/ins m1_n8607_n8040# out pass1u05u$3_1/ins
+ vss nfet$408
Xinv1u05u$3_0 vdd s4 vss inv1u05u$3_0/out inv1u05u$3
Xpass1u05u$3_4 vdd vss pass1u05u$3_7/ind pass1u05u$3_4/ins s2 inv1u05u$3_2/out pass1u05u$3
Xnfet$407_3 down down vss vss m1_n8807_n11192# vss nfet$407
Xpfet$381_15 m1_n8156_628# m1_n8156_628# pass1u05u$3_7/ins out out vdd pass1u05u$3_7/ins
+ m1_n8156_628# pass1u05u$3_7/ins pass1u05u$3_7/ins m1_n8156_628# out pass1u05u$3_7/ins
+ pass1u05u$3_7/ins pfet$381
Xnfet$408_15 vss down vss m1_n8607_n8040# down vss nfet$408
Xinv1u05u$3_1 vdd s3 vss inv1u05u$3_1/out inv1u05u$3
Xpass1u05u$3_5 vdd vss pass1u05u$3_7/ind pass1u05u$3_5/ins s3 inv1u05u$3_1/out pass1u05u$3
Xnfet$407_4 vss vss vss vss vss vss nfet$407
Xpfet$381_16 m1_n8156_628# m1_n8156_628# pass1u05u$3_7/ins out out vdd pass1u05u$3_7/ins
+ m1_n8156_628# pass1u05u$3_7/ins pass1u05u$3_7/ins m1_n8156_628# out pass1u05u$3_7/ins
+ pass1u05u$3_7/ins pfet$381
.ends

.subckt nfet$453 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$427 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$425 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$418 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$430 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$456 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$423 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt nfet$449 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$454 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt pfet$421 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$447 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$452 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$445 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$450 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$443 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$428 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt pfet$426 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt pfet$419 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$424 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$455 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt pfet$422 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$448 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt pfet$420 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$446 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$451 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt nfet$444 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$429 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt asc_PFD_DFF_20250831$2 vss down up vdd fdiv fref
Xnfet$453_9 m1_n5427_n10882# vss m1_n3884_n11124# vss nfet$453
Xpfet$427_2 vdd m1_1095_n11125# m1_832_n8573# m1_n3884_n11124# pfet$427
Xpfet$427_3 vdd m1_1452_n8889# m1_2556_n10129# m1_n3884_n9085# pfet$427
Xpfet$425_0 vdd m1_n5428_n3533# vdd m1_n5650_n4045# pfet$425
Xpfet$427_4 vdd vdd m1_1452_n8889# m1_832_n8573# pfet$427
Xpfet$418_0 vdd m1_832_n5785# m1_1096_n5165# m1_n3885_n6084# pfet$418
Xpfet$425_1 vdd vdd m1_n5428_n3533# m1_n4678_n3849# pfet$425
Xpfet$427_5 vdd vdd m1_1095_n11125# vdd pfet$427
Xpfet$418_1 vdd m1_1452_n5483# m1_2556_n4049# m1_n3885_n6084# pfet$418
Xpfet$430_0 vdd m1_5895_n8089# vdd down pfet$430
Xpfet$425_2 vdd m1_n5428_n5842# vdd m1_n5868_n3849# pfet$425
Xpfet$427_6 vdd vdd m1_1096_n9089# m1_1452_n8889# pfet$427
Xnfet$456_0 up up m1_5895_n8089# m1_5895_n8089# m1_5043_n9245# vss nfet$456
Xpfet$418_2 vdd m1_1095_n4045# m1_832_n5785# m1_n3885_n4045# pfet$418
Xpfet$425_3 vdd vdd m1_n5428_n5842# m1_n4678_n5482# pfet$425
Xpfet$430_1 vdd vdd m1_5895_n8089# up pfet$430
Xpfet$423_0 m1_n1926_n4095# vdd vdd m1_n3099_n4095# pfet$423
Xnfet$456_1 down down vss vss m1_5043_n9245# vss nfet$456
Xnfet$449_0 m1_n5428_n3533# vss m1_n3885_n4045# vss nfet$449
Xpfet$427_7 vdd m1_832_n8573# m1_1096_n9089# m1_n3884_n9085# pfet$427
Xpfet$418_3 vdd m1_2556_n4049# m1_3349_n5165# m1_n3885_n4045# pfet$418
Xpfet$423_1 m1_n4678_n3849# vdd vdd m1_n1926_n5680# pfet$423
Xnfet$449_1 m1_n5868_n3849# vss m1_n5650_n4045# vss nfet$449
Xpfet$427_8 vdd m1_1096_n9089# vdd m1_2068_n8889# pfet$427
Xpfet$423_2 m1_n1926_n5680# vdd vdd m1_n3099_n5680# pfet$423
Xnfet$449_2 m1_n5428_n5842# vss m1_n3885_n6084# vss nfet$449
Xpfet$427_9 vdd vdd m1_2068_n8889# m1_2758_n8889# pfet$427
Xnfet$454_0 m1_n3884_n11124# vss m1_n3098_n10720# vss nfet$454
Xpfet$423_3 m1_n4678_n5482# vdd vdd m1_n1926_n4095# pfet$423
Xpfet$421_0 vdd vdd m1_2758_n8889# m1_4978_n5483# pfet$421
Xnfet$449_3 fref vss m1_n5868_n3849# vss nfet$449
Xnfet$454_1 m1_n3884_n9085# vss m1_n3098_n9135# vss nfet$454
Xnfet$447_0 m1_5895_n8089# vss m1_5464_n5483# vss nfet$447
Xnfet$447_1 m1_5464_n5483# vss m1_4978_n5483# vss nfet$447
Xnfet$452_0 m1_2556_n10129# m1_2556_n10129# vss vss m1_3015_n10205# vss nfet$452
Xnfet$452_1 m1_1452_n8889# m1_1452_n8889# m1_1096_n9089# m1_1096_n9089# m1_1550_n9245#
+ vss nfet$452
Xnfet$445_0 m1_2779_n3533# vss up vss nfet$445
Xnfet$452_2 m1_2068_n8889# m1_2068_n8889# vss vss m1_1550_n9245# vss nfet$452
Xnfet$445_1 m1_2779_n3533# vss m1_3349_n5165# vss nfet$445
Xpfet$427_20 vdd m1_n5427_n8573# vdd m1_n5867_n10544# pfet$427
Xnfet$445_2 m1_2758_n8889# vss m1_2068_n5361# vss nfet$445
Xnfet$452_3 m1_2068_n8889# m1_2068_n8889# m1_2779_n10883# m1_2779_n10883# m1_3015_n10205#
+ vss nfet$452
Xnfet$450_0 m1_n4678_n3849# m1_n4678_n3849# m1_n5428_n3533# m1_n5428_n3533# m1_n5192_n4205#
+ vss nfet$450
Xpfet$427_10 vdd vdd m1_3349_n9089# m1_2779_n10883# pfet$427
Xnfet$445_3 m1_832_n5785# vss m1_1452_n5483# vss nfet$445
Xnfet$443_0 m1_n3885_n4045# m1_832_n5785# m1_1096_n5165# vss nfet$443
Xnfet$452_4 m1_n4677_n10522# m1_n4677_n10522# m1_n5427_n10882# m1_n5427_n10882# m1_n5191_n10204#
+ vss nfet$452
Xpfet$428_0 vdd vdd m1_n3098_n10720# m1_n3884_n11124# pfet$428
Xnfet$450_1 m1_n5650_n4045# m1_n5650_n4045# vss vss m1_n5192_n4205# vss nfet$450
Xpfet$427_11 vdd vdd down m1_2779_n10883# pfet$427
Xnfet$445_4 vdd vss m1_1095_n4045# vss nfet$445
Xnfet$452_5 m1_n5649_n11124# m1_n5649_n11124# vss vss m1_n5191_n10204# vss nfet$452
Xnfet$443_1 m1_n3885_n4045# m1_1452_n5483# m1_2556_n4049# vss nfet$443
Xpfet$428_1 vdd vdd m1_n3098_n9135# m1_n3884_n9085# pfet$428
Xnfet$450_2 m1_n4678_n5482# m1_n4678_n5482# m1_n5428_n5842# m1_n5428_n5842# m1_n5192_n5164#
+ vss nfet$450
Xpfet$427_12 vdd m1_2556_n10129# m1_3349_n9089# m1_n3884_n11124# pfet$427
Xnfet$443_2 m1_n3885_n6084# m1_1095_n4045# m1_832_n5785# vss nfet$443
Xnfet$452_6 m1_n4677_n8889# m1_n4677_n8889# m1_n5427_n8573# m1_n5427_n8573# m1_n5191_n9245#
+ vss nfet$452
Xnfet$450_3 m1_n5868_n3849# m1_n5868_n3849# vss vss m1_n5192_n5164# vss nfet$450
Xpfet$427_13 vdd vdd m1_n5427_n8573# m1_n4677_n8889# pfet$427
Xnfet$452_7 m1_n5867_n10544# m1_n5867_n10544# vss vss m1_n5191_n9245# vss nfet$452
Xnfet$443_3 m1_n3885_n6084# m1_2556_n4049# m1_3349_n5165# vss nfet$443
Xpfet$427_14 vdd vdd m1_n3884_n11124# m1_n5427_n10882# pfet$427
Xpfet$426_0 vdd vdd m1_n3099_n4095# m1_n3885_n4045# pfet$426
Xpfet$419_0 vdd vdd m1_1096_n5165# m1_1452_n5483# pfet$419
Xpfet$426_1 vdd vdd m1_n3099_n5680# m1_n3885_n6084# pfet$426
Xpfet$427_15 vdd m1_n5427_n10882# vdd m1_n5649_n11124# pfet$427
Xpfet$419_1 vdd m1_1096_n5165# vdd m1_2068_n5361# pfet$419
Xpfet$427_16 vdd vdd m1_n5427_n10882# m1_n4677_n10522# pfet$427
Xpfet$419_2 vdd m1_2779_n3533# vdd m1_2556_n4049# pfet$419
Xpfet$427_17 vdd vdd m1_n5649_n11124# m1_n5867_n10544# pfet$427
Xpfet$424_0 vdd vdd m1_n3885_n4045# m1_n5428_n3533# pfet$424
Xnfet$453_10 m1_n5867_n10544# vss m1_n5649_n11124# vss nfet$453
Xpfet$419_3 vdd vdd m1_2779_n3533# m1_2068_n5361# pfet$419
Xpfet$427_18 vdd vdd m1_n5867_n10544# fdiv pfet$427
Xpfet$424_1 vdd vdd m1_n5650_n4045# m1_n5868_n3849# pfet$424
Xnfet$453_11 fdiv vss m1_n5867_n10544# vss nfet$453
Xpfet$427_19 vdd vdd m1_n3884_n9085# m1_n5427_n8573# pfet$427
Xpfet$424_2 vdd vdd m1_n3885_n6084# m1_n5428_n5842# pfet$424
Xnfet$455_0 m1_n4677_n8889# m1_n1925_n10720# vss vss nfet$455
Xnfet$453_12 m1_n5427_n8573# vss m1_n3884_n9085# vss nfet$453
Xpfet$424_3 vdd vdd m1_n5868_n3849# fref pfet$424
Xpfet$422_0 vdd vdd m1_5464_n5483# m1_5895_n8089# pfet$422
Xnfet$455_1 m1_n1925_n10720# m1_n3098_n10720# vss vss nfet$455
Xnfet$448_0 m1_n1926_n4095# m1_n3099_n4095# vss vss nfet$448
Xpfet$422_1 vdd vdd m1_4978_n5483# m1_5464_n5483# pfet$422
Xnfet$455_2 m1_n4677_n10522# m1_n1925_n9135# vss vss nfet$455
Xnfet$448_1 m1_n4678_n3849# m1_n1926_n5680# vss vss nfet$448
Xnfet$455_3 m1_n1925_n9135# m1_n3098_n9135# vss vss nfet$455
Xnfet$448_2 m1_n1926_n5680# m1_n3099_n5680# vss vss nfet$448
Xnfet$453_0 m1_n3884_n9085# m1_1095_n11125# m1_832_n8573# vss nfet$453
Xpfet$420_0 vdd vdd m1_3349_n5165# m1_2779_n3533# pfet$420
Xnfet$453_1 m1_n3884_n11124# m1_1452_n8889# m1_2556_n10129# vss nfet$453
Xnfet$448_3 m1_n4678_n5482# m1_n1926_n4095# vss vss nfet$448
Xnfet$446_0 m1_4978_n5483# vss m1_2758_n8889# vss nfet$446
Xpfet$420_1 vdd vdd up m1_2779_n3533# pfet$420
Xnfet$453_2 m1_832_n8573# vss m1_1452_n8889# vss nfet$453
Xpfet$420_2 vdd vdd m1_2068_n5361# m1_2758_n8889# pfet$420
Xnfet$453_3 vdd vss m1_1095_n11125# vss nfet$453
Xnfet$451_0 m1_n3885_n4045# vss m1_n3099_n4095# vss nfet$451
Xpfet$420_3 vdd vdd m1_1452_n5483# m1_832_n5785# pfet$420
Xnfet$453_4 m1_n3884_n11124# m1_832_n8573# m1_1096_n9089# vss nfet$453
Xnfet$444_0 m1_2068_n5361# m1_2068_n5361# vss vss m1_1550_n5165# vss nfet$444
Xpfet$429_0 m1_n4677_n8889# vdd vdd m1_n1925_n10720# pfet$429
Xnfet$451_1 m1_n3885_n6084# vss m1_n3099_n5680# vss nfet$451
Xpfet$420_4 vdd vdd m1_1095_n4045# vdd pfet$420
Xnfet$453_5 m1_2758_n8889# vss m1_2068_n8889# vss nfet$453
Xnfet$444_1 m1_1452_n5483# m1_1452_n5483# m1_1096_n5165# m1_1096_n5165# m1_1550_n5165#
+ vss nfet$444
Xpfet$429_1 m1_n1925_n10720# vdd vdd m1_n3098_n10720# pfet$429
Xnfet$453_6 m1_2779_n10883# vss down vss nfet$453
Xnfet$444_2 m1_2556_n4049# m1_2556_n4049# vss vss m1_3015_n4205# vss nfet$444
Xpfet$429_2 m1_n4677_n10522# vdd vdd m1_n1925_n9135# pfet$429
Xnfet$444_3 m1_2068_n5361# m1_2068_n5361# m1_2779_n3533# m1_2779_n3533# m1_3015_n4205#
+ vss nfet$444
Xnfet$453_7 m1_2779_n10883# vss m1_3349_n9089# vss nfet$453
Xpfet$429_3 m1_n1925_n9135# vdd vdd m1_n3098_n9135# pfet$429
Xpfet$427_0 vdd vdd m1_2779_n10883# m1_2068_n8889# pfet$427
Xnfet$453_8 m1_n3884_n9085# m1_2556_n10129# m1_3349_n9089# vss nfet$453
Xpfet$427_1 vdd m1_2779_n10883# vdd m1_2556_n10129# pfet$427
.ends

.subckt pfet$409 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$412 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$438 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$410 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$436 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt nfet$434 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$413 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$411 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$437 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$435 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt asc_drive_buffer_up$2 vss out in vdd
Xpfet$409_0 out out m1_778_712# vdd m1_778_712# out vdd vdd m1_778_712# out m1_778_712#
+ m1_778_712# out m1_778_712# vdd m1_778_712# vdd m1_778_712# pfet$409
Xpfet$412_0 vdd vdd m1_n30_1318# m1_n566_1318# pfet$412
Xnfet$438_0 in vss m1_n566_1318# vss nfet$438
Xpfet$410_0 m1_778_712# vdd vdd m1_778_712# m1_506_712# m1_506_712# m1_778_712# vdd
+ m1_506_712# m1_506_712# pfet$410
Xnfet$436_0 m1_n30_1318# vss m1_506_712# vss nfet$436
Xnfet$434_0 m1_778_712# vss m1_506_712# m1_506_712# m1_506_712# m1_778_712# m1_778_712#
+ vss m1_506_712# vss nfet$434
Xpfet$413_0 vdd vdd m1_n566_1318# in pfet$413
Xpfet$411_0 vdd vdd m1_506_712# m1_n30_1318# pfet$411
Xnfet$437_0 m1_n566_1318# vss m1_n30_1318# vss nfet$437
Xnfet$435_0 out out vss m1_778_712# m1_778_712# out vss m1_778_712# m1_778_712# m1_778_712#
+ out m1_778_712# m1_778_712# out vss m1_778_712# vss vss nfet$435
.ends

.subckt pfet$431 a_254_0# a_348_560# w_n180_n88# a_414_0# a_n92_0# a_94_0# a_574_0#
+ a_508_560# a_188_560# a_28_560#
X0 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$457 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt BIAS$2 vdd vss 100n 200n res 200p1 200p2
Xpfet$431_10 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$431
Xpfet$431_11 vdd res vdd 200n vdd 200n vdd res res res pfet$431
Xpfet$431_12 vdd res vdd 100n vdd 100n vdd res res res pfet$431
Xpfet$431_13 vdd res vdd res vdd res vdd res res res pfet$431
Xpfet$431_14 vdd res vdd 200n vdd 200n vdd res res res pfet$431
Xpfet$431_15 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$431
Xpfet$431_0 vdd res vdd 200n vdd 200n vdd res res res pfet$431
Xnfet$457_0 m1_27_n1423# vss 200p1 m1_27_n1423# vss 200p1 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$457
Xpfet$431_1 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$431
Xnfet$457_1 vss vss vss vss vss vss vss vss vss vss nfet$457
Xpfet$431_3 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$431
Xpfet$431_2 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$431
Xnfet$457_2 m1_27_n1423# vss 200p2 m1_27_n1423# vss 200p2 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$457
Xpfet$431_4 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$431
Xnfet$457_3 vss vss vss vss vss vss vss vss vss vss nfet$457
Xpfet$431_5 vdd res vdd 200n vdd 200n vdd res res res pfet$431
Xnfet$457_4 m1_27_n1423# vss 200p2 m1_27_n1423# vss 200p2 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$457
Xnfet$457_6 m1_27_n1423# vss m1_27_n1423# m1_27_n1423# vss m1_27_n1423# m1_27_n1423#
+ vss m1_27_n1423# vss nfet$457
Xpfet$431_6 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$431
Xnfet$457_5 m1_27_n1423# vss 200p1 m1_27_n1423# vss 200p1 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$457
Xnfet$457_7 m1_27_n1423# vss m1_27_n1423# m1_27_n1423# vss m1_27_n1423# m1_27_n1423#
+ vss m1_27_n1423# vss nfet$457
Xpfet$431_7 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$431
Xpfet$431_8 vdd res vdd res vdd res vdd res res res pfet$431
Xpfet$431_9 vdd res vdd 100n vdd 100n vdd res res res pfet$431
.ends

.subckt pfet$402 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$393 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$428 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$400 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$398 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$426 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$419 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$431 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$396 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$424 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$417 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$422 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$394 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$420 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$392 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$405 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$403 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$429 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$401 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$399 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$427 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$425 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$397 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$418 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt nfet$430 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$423 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$395 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$421 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$406 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$404 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt asc_lock_detector_20250826$2 ref vdd div vss lock
Xpfet$402_0 vdd vdd m1_n8022_5099# m1_n10260_7868# pfet$402
Xpfet$393_7 vdd vdd m1_11370_4493# m1_10834_5099# pfet$393
Xnfet$428_0 div m1_n4030_5270# vss vss nfet$428
Xpfet$402_1 vdd vdd m1_n16410_5099# div pfet$402
Xnfet$428_1 m1_n6066_7868# vss m1_n4030_5270# vss nfet$428
Xpfet$402_2 vdd vdd m1_n12216_5099# m1_n14454_7868# pfet$402
Xpfet$400_0 m1_n11408_4493# vdd vdd m1_n11408_4493# m1_n11680_4493# m1_n11680_4493#
+ m1_n11408_4493# vdd m1_n11680_4493# m1_n11680_4493# pfet$400
Xpfet$398_0 vdd m1_17926_34# vdd m1_17703_788# pfet$398
Xnfet$426_0 m1_15979_2344# vss m1_16599_2028# vss nfet$426
Xpfet$400_1 m1_n7214_4493# vdd vdd m1_n7214_4493# m1_n7486_4493# m1_n7486_4493# m1_n7214_4493#
+ vdd m1_n7486_4493# m1_n7486_4493# pfet$400
Xpfet$398_1 vdd vdd m1_17926_34# m1_17215_2028# pfet$398
Xnfet$426_1 m1_15618_394# vss m1_15755_n208# vss nfet$426
Xnfet$419_0 m1_3254_n340# vss m1_2982_n340# m1_2982_n340# m1_2982_n340# m1_3254_n340#
+ m1_3254_n340# vss m1_2982_n340# vss nfet$419
Xpfet$400_2 m1_n15602_4493# vdd vdd m1_n15602_4493# m1_n15874_4493# m1_n15874_4493#
+ m1_n15602_4493# vdd m1_n15874_4493# m1_n15874_4493# pfet$400
Xnfet$426_2 m1_n2336_5099# vss m1_16242_n208# vss nfet$426
Xnfet$419_1 m1_7448_n340# vss m1_7176_n340# m1_7176_n340# m1_7176_n340# m1_7448_n340#
+ m1_7448_n340# vss m1_7176_n340# vss nfet$419
Xpfet$398_2 vdd m1_16243_1828# vdd m1_17215_2028# pfet$398
Xnfet$431_0 m1_19675_2344# vss lock vss nfet$431
Xpfet$396_0 vdd vdd m1_16599_2028# m1_15979_2344# pfet$396
Xpfet$398_3 vdd vdd m1_16243_1828# m1_16599_2028# pfet$398
Xnfet$426_3 m1_17926_34# vss m1_18496_1828# vss nfet$426
Xnfet$419_2 m1_11642_n340# vss m1_11370_n340# m1_11370_n340# m1_11370_n340# m1_11642_n340#
+ m1_11642_n340# vss m1_11370_n340# vss nfet$419
Xnfet$424_0 m1_15755_n208# m1_16599_2028# m1_17703_788# vss nfet$424
Xpfet$398_4 vdd m1_16243_5840# vdd m1_17215_5644# pfet$398
Xpfet$396_10 vdd vdd m1_15618_7156# m1_12790_7868# pfet$396
Xpfet$396_1 vdd vdd m1_16242_n208# m1_n2336_5099# pfet$396
Xnfet$424_1 m1_15618_394# m1_16242_n208# m1_15979_2344# vss nfet$424
Xnfet$417_0 m1_8596_n340# m1_8596_n340# vss m1_7448_n340# m1_7448_n340# m1_8596_n340#
+ vss m1_7448_n340# m1_7448_n340# m1_7448_n340# m1_8596_n340# m1_7448_n340# m1_7448_n340#
+ m1_8596_n340# vss m1_7448_n340# vss vss nfet$417
Xnfet$426_4 m1_12790_n340# vss m1_15618_394# vss nfet$426
Xnfet$419_3 m1_n940_n340# vss m1_n1212_n340# m1_n1212_n340# m1_n1212_n340# m1_n940_n340#
+ m1_n940_n340# vss m1_n1212_n340# vss nfet$419
Xnfet$419_4 m1_11642_4493# vss m1_11370_4493# m1_11370_4493# m1_11370_4493# m1_11642_4493#
+ m1_11642_4493# vss m1_11370_4493# vss nfet$419
Xpfet$398_5 vdd vdd m1_16243_5840# m1_16599_5522# pfet$398
Xpfet$396_2 vdd vdd m1_15755_n208# m1_15618_394# pfet$396
Xnfet$426_5 vss vss m1_17215_2028# vss nfet$426
Xpfet$396_11 vdd vdd m1_16599_5522# m1_15979_5220# pfet$396
Xnfet$417_1 m1_4402_n340# m1_4402_n340# vss m1_3254_n340# m1_3254_n340# m1_4402_n340#
+ vss m1_3254_n340# m1_3254_n340# m1_3254_n340# m1_4402_n340# m1_3254_n340# m1_3254_n340#
+ m1_4402_n340# vss m1_3254_n340# vss vss nfet$417
Xnfet$424_2 m1_15618_394# m1_17703_788# m1_18496_1828# vss nfet$424
Xpfet$398_6 vdd m1_17926_7472# vdd m1_17703_6956# pfet$398
Xnfet$419_5 m1_7448_4493# vss m1_7176_4493# m1_7176_4493# m1_7176_4493# m1_7448_4493#
+ m1_7448_4493# vss m1_7176_4493# vss nfet$419
Xpfet$396_12 vdd vdd m1_16242_6960# ref pfet$396
Xpfet$396_3 vdd vdd m1_18496_1828# m1_17926_34# pfet$396
Xnfet$417_2 m1_12790_n340# m1_12790_n340# vss m1_11642_n340# m1_11642_n340# m1_12790_n340#
+ vss m1_11642_n340# m1_11642_n340# m1_11642_n340# m1_12790_n340# m1_11642_n340# m1_11642_n340#
+ m1_12790_n340# vss m1_11642_n340# vss vss nfet$417
Xnfet$424_3 m1_15755_n208# m1_15979_2344# m1_16243_1828# vss nfet$424
Xnfet$426_6 m1_17926_34# vss m1_19469_1832# vss nfet$426
Xnfet$422_0 m1_n7214_4493# vss m1_n7486_4493# m1_n7486_4493# m1_n7486_4493# m1_n7214_4493#
+ m1_n7214_4493# vss m1_n7486_4493# vss nfet$422
Xpfet$394_0 m1_8596_n340# m1_8596_n340# m1_7448_n340# vdd m1_7448_n340# m1_8596_n340#
+ vdd vdd m1_7448_n340# m1_8596_n340# m1_7448_n340# m1_7448_n340# m1_8596_n340# m1_7448_n340#
+ vdd m1_7448_n340# vdd m1_7448_n340# pfet$394
Xnfet$419_6 m1_n940_4493# vss m1_n1212_4493# m1_n1212_4493# m1_n1212_4493# m1_n940_4493#
+ m1_n940_4493# vss m1_n1212_4493# vss nfet$419
Xpfet$398_7 vdd vdd m1_17926_7472# m1_17215_5644# pfet$398
Xpfet$396_4 vdd vdd m1_15618_394# m1_12790_n340# pfet$396
Xnfet$426_7 vss vss m1_17215_5644# vss nfet$426
Xpfet$396_13 vdd vdd m1_15755_6960# m1_15618_7156# pfet$396
Xnfet$424_4 m1_15618_7156# m1_17703_6956# m1_18496_5840# vss nfet$424
Xpfet$394_1 m1_12790_n340# m1_12790_n340# m1_11642_n340# vdd m1_11642_n340# m1_12790_n340#
+ vdd vdd m1_11642_n340# m1_12790_n340# m1_11642_n340# m1_11642_n340# m1_12790_n340#
+ m1_11642_n340# vdd m1_11642_n340# vdd m1_11642_n340# pfet$394
Xnfet$417_3 m1_208_n340# m1_208_n340# vss m1_n940_n340# m1_n940_n340# m1_208_n340#
+ vss m1_n940_n340# m1_n940_n340# m1_n940_n340# m1_208_n340# m1_n940_n340# m1_n940_n340#
+ m1_208_n340# vss m1_n940_n340# vss vss nfet$417
Xnfet$422_1 m1_n15602_4493# vss m1_n15874_4493# m1_n15874_4493# m1_n15874_4493# m1_n15602_4493#
+ m1_n15602_4493# vss m1_n15874_4493# vss nfet$422
Xnfet$419_7 m1_3254_4493# vss m1_2982_4493# m1_2982_4493# m1_2982_4493# m1_3254_4493#
+ m1_3254_4493# vss m1_2982_4493# vss nfet$419
Xnfet$417_4 m1_12790_7868# m1_12790_7868# vss m1_11642_4493# m1_11642_4493# m1_12790_7868#
+ vss m1_11642_4493# m1_11642_4493# m1_11642_4493# m1_12790_7868# m1_11642_4493# m1_11642_4493#
+ m1_12790_7868# vss m1_11642_4493# vss vss nfet$417
Xnfet$424_5 m1_15755_6960# m1_15979_5220# m1_16243_5840# vss nfet$424
Xnfet$426_8 m1_17926_7472# vss m1_19469_4920# vss nfet$426
Xpfet$396_5 vdd vdd m1_17215_2028# vss pfet$396
Xnfet$422_2 m1_n11408_4493# vss m1_n11680_4493# m1_n11680_4493# m1_n11680_4493# m1_n11408_4493#
+ m1_n11408_4493# vss m1_n11680_4493# vss nfet$422
Xpfet$394_2 m1_4402_n340# m1_4402_n340# m1_3254_n340# vdd m1_3254_n340# m1_4402_n340#
+ vdd vdd m1_3254_n340# m1_4402_n340# m1_3254_n340# m1_3254_n340# m1_4402_n340# m1_3254_n340#
+ vdd m1_3254_n340# vdd m1_3254_n340# pfet$394
Xnfet$426_9 m1_17926_7472# vss m1_18496_5840# vss nfet$426
Xnfet$417_5 m1_8596_7868# m1_8596_7868# vss m1_7448_4493# m1_7448_4493# m1_8596_7868#
+ vss m1_7448_4493# m1_7448_4493# m1_7448_4493# m1_8596_7868# m1_7448_4493# m1_7448_4493#
+ m1_8596_7868# vss m1_7448_4493# vss vss nfet$417
Xnfet$424_6 m1_15618_7156# m1_16242_6960# m1_15979_5220# vss nfet$424
Xpfet$396_6 vdd vdd m1_19469_1832# m1_17926_34# pfet$396
Xpfet$394_3 m1_208_n340# m1_208_n340# m1_n940_n340# vdd m1_n940_n340# m1_208_n340#
+ vdd vdd m1_n940_n340# m1_208_n340# m1_n940_n340# m1_n940_n340# m1_208_n340# m1_n940_n340#
+ vdd m1_n940_n340# vdd m1_n940_n340# pfet$394
Xnfet$420_0 m1_n6066_7868# m1_n6066_7868# vss m1_n7214_4493# m1_n7214_4493# m1_n6066_7868#
+ vss m1_n7214_4493# m1_n7214_4493# m1_n7214_4493# m1_n6066_7868# m1_n7214_4493# m1_n7214_4493#
+ m1_n6066_7868# vss m1_n7214_4493# vss vss nfet$420
Xpfet$392_0 vdd vdd m1_6640_1478# m1_4402_n340# pfet$392
Xpfet$405_0 vdd m1_19675_2344# vdd m1_19469_1832# pfet$405
Xpfet$396_7 vdd vdd m1_17215_5644# vss pfet$396
Xnfet$417_6 m1_208_7868# m1_208_7868# vss m1_n940_4493# m1_n940_4493# m1_208_7868#
+ vss m1_n940_4493# m1_n940_4493# m1_n940_4493# m1_208_7868# m1_n940_4493# m1_n940_4493#
+ m1_208_7868# vss m1_n940_4493# vss vss nfet$417
Xnfet$424_7 m1_15755_6960# m1_16599_5522# m1_17703_6956# vss nfet$424
Xpfet$392_1 vdd vdd m1_10834_1478# m1_8596_n340# pfet$392
Xpfet$394_4 m1_208_7868# m1_208_7868# m1_n940_4493# vdd m1_n940_4493# m1_208_7868#
+ vdd vdd m1_n940_4493# m1_208_7868# m1_n940_4493# m1_n940_4493# m1_208_7868# m1_n940_4493#
+ vdd m1_n940_4493# vdd m1_n940_4493# pfet$394
Xnfet$420_1 m1_n14454_7868# m1_n14454_7868# vss m1_n15602_4493# m1_n15602_4493# m1_n14454_7868#
+ vss m1_n15602_4493# m1_n15602_4493# m1_n15602_4493# m1_n14454_7868# m1_n15602_4493#
+ m1_n15602_4493# m1_n14454_7868# vss m1_n15602_4493# vss vss nfet$420
Xpfet$405_1 vdd vdd m1_19675_2344# m1_19469_4920# pfet$405
Xnfet$417_7 m1_4402_7868# m1_4402_7868# vss m1_3254_4493# m1_3254_4493# m1_4402_7868#
+ vss m1_3254_4493# m1_3254_4493# m1_3254_4493# m1_4402_7868# m1_3254_4493# m1_3254_4493#
+ m1_4402_7868# vss m1_3254_4493# vss vss nfet$417
Xpfet$394_5 m1_12790_7868# m1_12790_7868# m1_11642_4493# vdd m1_11642_4493# m1_12790_7868#
+ vdd vdd m1_11642_4493# m1_12790_7868# m1_11642_4493# m1_11642_4493# m1_12790_7868#
+ m1_11642_4493# vdd m1_11642_4493# vdd m1_11642_4493# pfet$394
Xpfet$396_8 vdd vdd m1_19469_4920# m1_17926_7472# pfet$396
Xnfet$420_2 m1_n10260_7868# m1_n10260_7868# vss m1_n11408_4493# m1_n11408_4493# m1_n10260_7868#
+ vss m1_n11408_4493# m1_n11408_4493# m1_n11408_4493# m1_n10260_7868# m1_n11408_4493#
+ m1_n11408_4493# m1_n10260_7868# vss m1_n11408_4493# vss vss nfet$420
Xpfet$392_2 vdd vdd m1_n1748_1478# ref pfet$392
Xpfet$396_9 vdd vdd m1_18496_5840# m1_17926_7472# pfet$396
Xpfet$394_6 m1_4402_7868# m1_4402_7868# m1_3254_4493# vdd m1_3254_4493# m1_4402_7868#
+ vdd vdd m1_3254_4493# m1_4402_7868# m1_3254_4493# m1_3254_4493# m1_4402_7868# m1_3254_4493#
+ vdd m1_3254_4493# vdd m1_3254_4493# pfet$394
Xpfet$392_3 vdd vdd m1_n1748_5099# m1_n2336_5099# pfet$392
Xpfet$403_0 vdd vdd vdd m1_n3798_6028# div div pfet$403
Xpfet$394_7 m1_8596_7868# m1_8596_7868# m1_7448_4493# vdd m1_7448_4493# m1_8596_7868#
+ vdd vdd m1_7448_4493# m1_8596_7868# m1_7448_4493# m1_7448_4493# m1_8596_7868# m1_7448_4493#
+ vdd m1_7448_4493# vdd m1_7448_4493# pfet$394
Xnfet$429_0 m1_n4030_5270# vss m1_n2336_5099# vss nfet$429
Xpfet$392_4 vdd vdd m1_6640_5099# m1_4402_7868# pfet$392
Xpfet$403_1 vdd m1_n4030_5270# m1_n4030_5270# m1_n3798_6028# m1_n6066_7868# m1_n6066_7868#
+ pfet$403
Xpfet$392_5 vdd vdd m1_10834_5099# m1_8596_7868# pfet$392
Xpfet$392_6 vdd vdd m1_2446_5099# m1_208_7868# pfet$392
Xnfet$426_10 m1_12790_7868# vss m1_15618_7156# vss nfet$426
Xpfet$401_0 vdd vdd m1_n11680_4493# m1_n12216_5099# pfet$401
Xpfet$399_0 m1_n10260_7868# m1_n10260_7868# m1_n11408_4493# vdd m1_n11408_4493# m1_n10260_7868#
+ vdd vdd m1_n11408_4493# m1_n10260_7868# m1_n11408_4493# m1_n11408_4493# m1_n10260_7868#
+ m1_n11408_4493# vdd m1_n11408_4493# vdd m1_n11408_4493# pfet$399
Xpfet$392_7 vdd vdd m1_2446_1478# m1_208_n340# pfet$392
Xnfet$427_0 m1_n14454_7868# vss m1_n12216_5099# vss nfet$427
Xnfet$426_11 m1_15979_5220# vss m1_16599_5522# vss nfet$426
Xpfet$401_1 vdd vdd m1_n7486_4493# m1_n8022_5099# pfet$401
Xnfet$427_1 div vss m1_n16410_5099# vss nfet$427
Xpfet$399_1 m1_n6066_7868# m1_n6066_7868# m1_n7214_4493# vdd m1_n7214_4493# m1_n6066_7868#
+ vdd vdd m1_n7214_4493# m1_n6066_7868# m1_n7214_4493# m1_n7214_4493# m1_n6066_7868#
+ m1_n7214_4493# vdd m1_n7214_4493# vdd m1_n7214_4493# pfet$399
Xnfet$426_12 m1_15618_7156# vss m1_15755_6960# vss nfet$426
Xpfet$401_2 vdd vdd m1_n15874_4493# m1_n16410_5099# pfet$401
Xpfet$399_2 m1_n14454_7868# m1_n14454_7868# m1_n15602_4493# vdd m1_n15602_4493# m1_n14454_7868#
+ vdd vdd m1_n15602_4493# m1_n14454_7868# m1_n15602_4493# m1_n15602_4493# m1_n14454_7868#
+ m1_n15602_4493# vdd m1_n15602_4493# vdd m1_n15602_4493# pfet$399
Xnfet$427_2 m1_n10260_7868# vss m1_n8022_5099# vss nfet$427
Xnfet$426_13 ref vss m1_16242_6960# vss nfet$426
Xnfet$425_0 m1_17215_2028# m1_17215_2028# m1_17926_34# m1_17926_34# m1_18162_712#
+ vss nfet$425
Xpfet$397_0 vdd m1_16599_2028# m1_17703_788# m1_15618_394# pfet$397
Xpfet$397_1 vdd m1_16242_n208# m1_15979_2344# m1_15755_n208# pfet$397
Xnfet$425_1 m1_17703_788# m1_17703_788# vss vss m1_18162_712# vss nfet$425
Xnfet$418_0 m1_10834_1478# vss m1_11370_n340# vss nfet$418
Xnfet$418_1 m1_2446_1478# vss m1_2982_n340# vss nfet$418
Xpfet$397_2 vdd m1_15979_2344# m1_16243_1828# m1_15618_394# pfet$397
Xnfet$425_2 m1_16599_2028# m1_16599_2028# m1_16243_1828# m1_16243_1828# m1_16697_1672#
+ vss nfet$425
Xnfet$430_0 m1_19469_4920# m1_19469_4920# m1_19675_2344# m1_19675_2344# m1_19911_1672#
+ vss nfet$430
Xpfet$397_3 vdd m1_17703_788# m1_18496_1828# m1_15755_n208# pfet$397
Xnfet$423_0 m1_8596_n340# vss m1_10834_1478# vss nfet$423
Xnfet$418_2 m1_6640_1478# vss m1_7176_n340# vss nfet$418
Xnfet$425_3 m1_17215_2028# m1_17215_2028# vss vss m1_16697_1672# vss nfet$425
Xpfet$395_0 m1_7448_n340# vdd vdd m1_7448_n340# m1_7176_n340# m1_7176_n340# m1_7448_n340#
+ vdd m1_7176_n340# m1_7176_n340# pfet$395
Xnfet$430_1 m1_19469_1832# m1_19469_1832# vss vss m1_19911_1672# vss nfet$430
Xpfet$397_4 vdd m1_17703_6956# m1_18496_5840# m1_15755_6960# pfet$397
Xpfet$395_1 m1_11642_n340# vdd vdd m1_11642_n340# m1_11370_n340# m1_11370_n340# m1_11642_n340#
+ vdd m1_11370_n340# m1_11370_n340# pfet$395
Xnfet$418_3 m1_n1748_1478# vss m1_n1212_n340# vss nfet$418
Xnfet$425_4 m1_17215_5644# m1_17215_5644# vss vss m1_16697_5840# vss nfet$425
Xnfet$423_1 m1_4402_n340# vss m1_6640_1478# vss nfet$423
Xpfet$397_5 vdd m1_15979_5220# m1_16243_5840# m1_15618_7156# pfet$397
Xnfet$418_4 m1_10834_5099# vss m1_11370_4493# vss nfet$418
Xnfet$425_5 m1_16599_5522# m1_16599_5522# m1_16243_5840# m1_16243_5840# m1_16697_5840#
+ vss nfet$425
Xpfet$395_2 m1_3254_n340# vdd vdd m1_3254_n340# m1_2982_n340# m1_2982_n340# m1_3254_n340#
+ vdd m1_2982_n340# m1_2982_n340# pfet$395
Xnfet$423_2 ref vss m1_n1748_1478# vss nfet$423
Xnfet$418_5 m1_6640_5099# vss m1_7176_4493# vss nfet$418
Xnfet$425_6 m1_17215_5644# m1_17215_5644# m1_17926_7472# m1_17926_7472# m1_18162_6800#
+ vss nfet$425
Xpfet$397_6 vdd m1_16599_5522# m1_17703_6956# m1_15618_7156# pfet$397
Xpfet$393_0 vdd vdd m1_7176_n340# m1_6640_1478# pfet$393
Xpfet$395_3 m1_n940_n340# vdd vdd m1_n940_n340# m1_n1212_n340# m1_n1212_n340# m1_n940_n340#
+ vdd m1_n1212_n340# m1_n1212_n340# pfet$395
Xnfet$423_3 m1_n2336_5099# vss m1_n1748_5099# vss nfet$423
Xnfet$421_0 m1_n8022_5099# vss m1_n7486_4493# vss nfet$421
Xpfet$406_0 vdd vdd lock m1_19675_2344# pfet$406
Xpfet$397_7 vdd m1_16242_6960# m1_15979_5220# m1_15755_6960# pfet$397
Xnfet$418_6 m1_n1748_5099# vss m1_n1212_4493# vss nfet$418
Xnfet$425_7 m1_17703_6956# m1_17703_6956# vss vss m1_18162_6800# vss nfet$425
Xpfet$395_4 m1_n940_4493# vdd vdd m1_n940_4493# m1_n1212_4493# m1_n1212_4493# m1_n940_4493#
+ vdd m1_n1212_4493# m1_n1212_4493# pfet$395
Xnfet$421_1 m1_n16410_5099# vss m1_n15874_4493# vss nfet$421
Xnfet$423_4 m1_8596_7868# vss m1_10834_5099# vss nfet$423
Xpfet$393_1 vdd vdd m1_11370_n340# m1_10834_1478# pfet$393
Xnfet$418_7 m1_2446_5099# vss m1_2982_4493# vss nfet$418
Xpfet$395_5 m1_11642_4493# vdd vdd m1_11642_4493# m1_11370_4493# m1_11370_4493# m1_11642_4493#
+ vdd m1_11370_4493# m1_11370_4493# pfet$395
Xnfet$423_5 m1_4402_7868# vss m1_6640_5099# vss nfet$423
Xpfet$393_2 vdd vdd m1_2982_n340# m1_2446_1478# pfet$393
Xnfet$421_2 m1_n12216_5099# vss m1_n11680_4493# vss nfet$421
Xpfet$395_6 m1_3254_4493# vdd vdd m1_3254_4493# m1_2982_4493# m1_2982_4493# m1_3254_4493#
+ vdd m1_2982_4493# m1_2982_4493# pfet$395
Xnfet$423_6 m1_208_n340# vss m1_2446_1478# vss nfet$423
Xpfet$393_3 vdd vdd m1_n1212_n340# m1_n1748_1478# pfet$393
Xpfet$404_0 vdd vdd m1_n2336_5099# m1_n4030_5270# pfet$404
Xnfet$423_7 m1_208_7868# vss m1_2446_5099# vss nfet$423
Xpfet$395_7 m1_7448_4493# vdd vdd m1_7448_4493# m1_7176_4493# m1_7176_4493# m1_7448_4493#
+ vdd m1_7176_4493# m1_7176_4493# pfet$395
Xpfet$393_4 vdd vdd m1_n1212_4493# m1_n1748_5099# pfet$393
Xpfet$393_5 vdd vdd m1_2982_4493# m1_2446_5099# pfet$393
Xpfet$393_6 vdd vdd m1_7176_4493# m1_6640_5099# pfet$393
.ends

.subckt pfet$389 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$387 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$415 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$413 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$390 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$388 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$416 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$414 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$391 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$412 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt asc_hysteresis_buffer$7 vss in vdd out
Xpfet$389_0 vdd vdd m1_348_648# in pfet$389
Xpfet$387_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd
+ m1_884_42# m1_884_42# pfet$387
Xnfet$415_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$415
Xnfet$413_0 m1_348_648# vss m1_884_42# vss nfet$413
Xpfet$390_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$390
Xpfet$388_0 vdd vdd m1_884_42# m1_348_648# pfet$388
Xnfet$416_0 m1_1156_42# vss m1_884_42# vss nfet$416
Xnfet$414_0 in vss m1_348_648# vss nfet$414
Xpfet$391_0 vdd vdd m1_884_42# m1_1156_42# pfet$391
Xnfet$412_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$412
.ends

.subckt pfet$432 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=9.75p pd=31.3u as=9.75p ps=31.3u w=15u l=0.5u
.ends

.subckt cap_mim$8 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
.ends

.subckt nfet$458 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.5u
.ends

.subckt nfet$459 a_n84_0# a_38_n132# a_138_0# VSUBS
X0 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.5u
.ends

.subckt pfet$433 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=9.75p pd=31.3u as=9.75p ps=31.3u w=15u l=0.5u
.ends

.subckt nfet$460 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$434 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt CSRVCO_20250823$2 vctrl vosc vdd vss
Xpfet$432_0 vdd vdd m1_n12264_2422# m1_n16019_266# pfet$432
Xcap_mim$8_3 vss m1_n11916_1270# cap_mim$8
Xnfet$458_0 m1_n9838_266# m1_n12754_674# m1_n9352_266# vss nfet$458
Xpfet$432_1 vdd vdd m1_n14208_3657# m1_n16019_266# pfet$432
Xcap_mim$8_4 vss m1_n9352_266# cap_mim$8
Xnfet$458_1 vctrl vss m1_n12268_985# vss nfet$458
Xpfet$432_2 vdd vdd m1_n13722_3340# m1_n16019_266# pfet$432
Xcap_mim$8_5 vss m1_n9838_266# cap_mim$8
Xnfet$458_3 vctrl vss m1_n13794_186# vss nfet$458
Xnfet$458_2 vctrl vss m1_n14283_186# vss nfet$458
Xcap_mim$8_6 vss m1_n11782_266# cap_mim$8
Xpfet$432_3 vdd m1_n16019_266# vdd m1_n16019_266# pfet$432
Xnfet$458_4 vctrl vss m1_n13240_368# vss nfet$458
Xpfet$432_4 vdd vdd m1_n13236_3035# m1_n16019_266# pfet$432
Xnfet$458_5 vctrl vss m1_n12754_674# vss nfet$458
Xpfet$432_5 vdd vdd m1_n14693_3963# m1_n16019_266# pfet$432
Xnfet$458_6 vctrl m1_n16019_266# vss vss nfet$458
Xpfet$432_6 vdd vdd m1_n12750_2729# m1_n16019_266# pfet$432
Xnfet$458_7 vctrl vss m1_n15245_186# vss nfet$458
Xpfet$432_8 vdd m1_n13236_3035# m1_n9838_266# m1_n10324_266# pfet$432
Xpfet$432_7 vdd vdd m1_n15180_4275# m1_n16019_266# pfet$432
Xnfet$458_8 vctrl vss m1_n14765_186# vss nfet$458
Xpfet$432_9 vdd m1_n12750_2729# m1_n9352_266# m1_n9838_266# pfet$432
Xnfet$458_10 m1_n9352_266# m1_n12268_985# m1_n11916_1270# vss nfet$458
Xnfet$458_9 m1_n10324_266# m1_n13240_368# m1_n9838_266# vss nfet$458
Xnfet$458_11 m1_n11916_1270# m1_n15245_186# m1_n11782_266# vss nfet$458
Xnfet$458_12 m1_n11782_266# m1_n14765_186# m1_n11296_266# vss nfet$458
Xnfet$458_13 m1_n11296_266# m1_n14283_186# m1_n10810_266# vss nfet$458
Xpfet$432_10 vdd m1_n14208_3657# m1_n10810_266# m1_n11296_266# pfet$432
Xnfet$458_14 m1_n10810_266# m1_n13794_186# m1_n10324_266# vss nfet$458
Xpfet$432_11 vdd m1_n12264_2422# m1_n11916_1270# m1_n9352_266# pfet$432
Xpfet$432_12 vdd m1_n14693_3963# m1_n11296_266# m1_n11782_266# pfet$432
Xnfet$459_0 vss vss vss vss nfet$459
Xpfet$432_13 vdd m1_n13722_3340# m1_n10324_266# m1_n10810_266# pfet$432
Xpfet$433_0 vdd vdd vdd vdd pfet$433
Xpfet$432_14 vdd m1_n15180_4275# m1_n11782_266# m1_n11916_1270# pfet$432
Xnfet$459_1 vss vss vss vss nfet$459
Xpfet$433_1 vdd vdd vdd vdd pfet$433
Xnfet$460_0 m1_n8380_274# vss vosc vss nfet$460
Xnfet$460_1 m1_n11916_1270# vss m1_n8380_274# vss nfet$460
Xpfet$434_1 vdd vdd m1_n8380_274# m1_n11916_1270# pfet$434
Xpfet$434_0 vdd vdd vosc m1_n8380_274# pfet$434
Xcap_mim$8_1 vss m1_n10810_266# cap_mim$8
Xcap_mim$8_0 vss m1_n11296_266# cap_mim$8
Xcap_mim$8_2 vss m1_n10324_266# cap_mim$8
.ends

.subckt xp_3_1_MUX$4 S0 S1 VDD VSS OUT_1 C_1 B_1 A_1
Xnfet$433_0 S1 VSS m1_n432_n1290# VSS nfet$433
Xnfet$433_1 S0 VSS m1_n432_458# VSS nfet$433
Xpfet$407_0 VDD A_1 m1_239_n318# m1_n432_458# pfet$407
Xpfet$407_2 VDD B_1 m1_239_n318# S0 pfet$407
Xpfet$407_1 VDD C_1 OUT_1 S1 pfet$407
Xpfet$407_3 VDD m1_239_n318# OUT_1 m1_n432_n1290# pfet$407
Xnfet$432_0 m1_n432_n1290# C_1 OUT_1 VSS nfet$432
Xnfet$432_1 m1_n432_458# B_1 m1_239_n318# VSS nfet$432
Xnfet$432_2 S1 m1_239_n318# OUT_1 VSS nfet$432
Xnfet$432_3 S0 A_1 m1_239_n318# VSS nfet$432
Xpfet$408_0 VDD VDD m1_n432_n1290# S1 pfet$408
Xpfet$408_1 VDD VDD m1_n432_458# S0 pfet$408
.ends

.subckt asc_dual_psd_def_20250809$4 vdd vss pd1 pd2 pd3 pd4 pd5 pd6 pd7 pd8 pd9 fout
+ sd1 sd2 sd3 sd4 sd5 sd6 sd7 sd8 sd9 fin define
Xpfet$356_6 vdd vdd m1_n290_24224# m1_n910_23922# pfet$356
Xpfet$349_5 vdd m1_7198_15778# m1_6377_16202# m1_6116_17343# pfet$349
Xnfet$371_6 m1_2384_21590# m1_2384_21590# m1_3871_22513# m1_3871_22513# m1_2843_21586#
+ vss nfet$371
Xnfet$378_10 m1_32675_25947# vss m1_35071_24542# vss nfet$378
Xpfet$351_19 vdd m1_n3822_20130# m1_n3822_20130# m1_27441_19850# m1_27003_19550# m1_27003_19550#
+ pfet$351
Xnfet$389_20 m1_22493_16080# m1_22493_16080# m1_22034_17714# m1_22034_17714# m1_22591_16398#
+ vss nfet$389
Xpfet$354_3 vdd vdd m1_5901_19550# m1_649_17714# pfet$354
Xnfet$375_11 m1_9331_15478# vss m1_15171_20152# vss nfet$375
Xpfet$352_0 vdd vdd m1_n1133_21590# m1_n1263_21786# pfet$352
Xnfet$389_7 m1_5761_16080# m1_5761_16080# m1_5302_17714# m1_5302_17714# m1_5859_16398#
+ vss nfet$389
Xnfet$396_8 m1_9624_19404# m1_9624_19404# vss vss m1_n3724_21430# vss nfet$396
Xpfet$349_108 vdd vdd m1_15454_18030# m1_15564_15778# pfet$349
Xnfet$372_12 m1_16452_19550# m1_16452_19550# vss vss m1_16890_20470# vss nfet$372
Xnfet$392_2 m1_n6274_17836# m1_n5351_15778# m1_n6172_16202# vss nfet$392
Xnfet$378_0 m1_n10452_25858# vss m1_n1271_25858# vss nfet$378
Xpfet$349_19 vdd m1_3015_15778# m1_2194_16202# m1_1933_17343# pfet$349
Xpfet$377_2 vdd m1_n5764_21786# m1_n5764_21786# m1_n5019_22344# m1_n5227_21418# m1_n5227_21418#
+ pfet$377
Xnfet$371_7 m1_5771_21786# m1_5771_21786# m1_7388_22513# m1_7388_22513# m1_6992_21586#
+ vss nfet$371
Xnfet$378_11 m1_32554_23922# vss m1_33174_24224# vss nfet$378
Xpfet$356_7 vdd vdd m1_32330_25662# m1_32193_25858# pfet$356
Xpfet$349_6 vdd vdd m1_7198_15778# m1_7555_16080# pfet$349
Xnfet$389_21 m1_14127_16080# m1_14127_16080# vss vss m1_15690_17358# vss nfet$389
Xnfet$389_10 m1_1578_16080# m1_1578_16080# m1_1119_17714# m1_1119_17714# m1_1676_16398#
+ vss nfet$389
Xpfet$354_4 vdd vdd m1_12935_19550# m1_9015_17714# pfet$354
Xnfet$375_12 m1_13514_15478# vss m1_18688_20152# vss nfet$375
Xpfet$352_1 vdd vdd m1_11671_21786# m1_11039_21786# pfet$352
Xnfet$389_8 m1_3015_15778# m1_3015_15778# m1_2905_18030# m1_2905_18030# m1_3141_17358#
+ vss nfet$389
Xnfet$396_9 m1_n6380_21786# m1_n6380_21786# m1_n6839_21786# m1_n6839_21786# m1_n6282_21430#
+ vss nfet$396
Xpfet$349_109 vdd vdd m1_10299_17343# m1_13198_17714# pfet$349
Xnfet$372_13 m1_19969_19550# m1_19969_19550# vss vss m1_20407_20470# vss nfet$372
Xnfet$397_10 vss vss m1_n4978_24224# vss nfet$397
Xnfet$392_3 m1_n6433_17343# m1_n6172_16202# m1_n6657_17518# vss nfet$392
Xnfet$378_1 m1_n789_25858# vss m1_n647_25662# vss nfet$378
Xnfet$371_8 m1_23486_21590# m1_23486_21590# m1_24973_22513# m1_24973_22513# m1_23945_21586#
+ vss nfet$371
Xnfet$378_12 m1_32675_25947# vss m1_28624_21786# vss nfet$378
Xpfet$356_8 vdd vdd m1_33174_24224# m1_32554_23922# pfet$356
Xnfet$390_0 m1_4620_20152# m1_4620_20152# m1_2590_19404# m1_2590_19404# m1_3454_20470#
+ vss nfet$390
Xpfet$349_7 vdd vdd m1_6275_17836# m1_6116_17343# pfet$349
Xpfet$375_0 vdd vdd m1_n7186_25858# m1_n10452_25858# pfet$375
Xpfet$354_5 vdd vdd m1_8137_20152# m1_965_15478# pfet$354
Xnfet$403_0 m1_n927_19404# m1_n927_19404# vss vss m1_n6282_20470# vss nfet$403
Xnfet$389_22 m1_15564_15778# m1_15564_15778# m1_15454_18030# m1_15454_18030# m1_15690_17358#
+ vss nfet$389
Xnfet$389_11 m1_6377_16202# m1_6377_16202# vss vss m1_5859_16398# vss nfet$389
Xnfet$375_13 m1_13198_17714# vss m1_16452_19550# vss nfet$375
Xpfet$352_2 vdd vdd m1_12935_21590# m1_12805_21786# pfet$352
Xnfet$389_9 m1_2194_16202# m1_2194_16202# vss vss m1_1676_16398# vss nfet$389
Xpfet$348_110 vdd m1_11903_24542# vdd m1_12875_24346# pfet$348
Xnfet$372_14 m1_17381_17714# m1_17381_17714# vss vss m1_21039_20470# vss nfet$372
Xnfet$397_11 m1_n10452_25858# vss m1_n4847_25662# vss nfet$397
Xnfet$392_4 m1_27031_17343# m1_27292_16202# m1_26807_17518# vss nfet$392
Xnfet$378_2 m1_n1271_25858# vss m1_n1134_25662# vss nfet$378
Xnfet$371_9 m1_23356_21786# m1_23356_21786# m1_24973_22513# m1_24973_22513# m1_24577_21586#
+ vss nfet$371
Xnfet$378_13 m1_32675_25947# vss m1_32817_25662# vss nfet$378
Xpfet$356_9 vdd vdd m1_28624_21786# m1_32675_25947# pfet$356
Xnfet$383_0 m1_21456_22513# m1_21456_22513# m1_30256_19792# m1_30256_19792# m1_30492_20470#
+ vss nfet$383
Xnfet$390_1 m1_1103_20152# m1_1103_20152# m1_n927_19404# m1_n927_19404# m1_n63_20470#
+ vss nfet$390
Xpfet$349_8 vdd vdd m1_9331_15478# sd5 pfet$349
Xpfet$368_0 vdd vdd m1_n7513_20152# m1_35837_22102# pfet$368
Xpfet$375_1 vdd m1_n7186_25858# vdd m1_n6111_25858# pfet$375
Xnfet$403_1 m1_n2543_20130# m1_n2543_20130# m1_n5227_20152# m1_n5227_20152# m1_n2445_20470#
+ vss nfet$403
Xnfet$389_23 m1_18926_16202# m1_18926_16202# vss vss m1_18408_16398# vss nfet$389
Xpfet$354_6 vdd vdd m1_9418_19550# m1_4832_17714# pfet$354
Xnfet$389_12 m1_n1168_15778# m1_n1168_15778# m1_n1278_18030# m1_n1278_18030# m1_n1042_17358#
+ vss nfet$389
Xnfet$370_80 m1_28147_25662# m1_28991_24224# m1_30095_25658# vss nfet$370
Xpfet$352_10 vdd vdd m1_23486_21590# m1_23356_21786# pfet$352
Xnfet$375_14 m1_21564_17714# vss m1_23486_19550# vss nfet$375
Xpfet$352_3 vdd vdd m1_9418_21590# m1_9288_21786# pfet$352
Xpfet$348_100 vdd vdd m1_29607_24346# m1_n7513_20152# pfet$348
Xpfet$350_0 vdd vdd vdd m1_n674_22102# m1_n1133_21590# m1_n1133_21590# pfet$350
Xnfet$372_15 m1_21564_17714# m1_21564_17714# vss vss m1_24556_20470# vss nfet$372
Xnfet$397_12 m1_n10452_25858# vss m1_n5571_25662# vss nfet$397
Xnfet$392_5 m1_27031_17343# m1_29087_15778# m1_28470_16080# vss nfet$392
Xnfet$378_3 m1_n7513_20152# vss m1_326_24346# vss nfet$378
Xnfet$373_80 m1_18824_17836# m1_19747_15778# m1_18926_16202# vss nfet$373
Xnfet$383_1 m1_14422_22513# m1_14422_22513# m1_31535_19792# m1_31535_19792# m1_31771_20470#
+ vss nfet$383
Xnfet$390_2 m1_n3218_15478# m1_n3218_15478# m1_2590_19404# m1_2590_19404# m1_2822_20470#
+ vss nfet$390
Xpfet$349_9 vdd vdd m1_8172_15778# m1_5302_17714# pfet$349
Xnfet$376_0 sd9 vss m1_n7401_15478# vss nfet$376
Xnfet$389_24 m1_18310_16080# m1_18310_16080# m1_17851_17714# m1_17851_17714# m1_18408_16398#
+ vss nfet$389
Xpfet$354_7 vdd vdd m1_11654_20152# m1_5148_15478# pfet$354
Xnfet$389_13 m1_n2605_16080# m1_n2605_16080# vss vss m1_n1042_17358# vss nfet$389
Xnfet$370_81 m1_n7513_20152# vss m1_25424_24346# vss nfet$370
Xnfet$370_70 m1_21590_21786# vss m1_28010_25858# vss nfet$370
Xpfet$352_11 vdd vdd m1_18705_21786# m1_18073_21786# pfet$352
Xpfet$380_0 vdd vdd m1_n8145_21908# m1_n6839_20152# pfet$380
Xnfet$375_15 m1_17697_15478# vss m1_22205_20152# vss nfet$375
Xpfet$352_4 vdd vdd m1_8154_21786# m1_7522_21786# pfet$352
Xpfet$350_1 vdd m1_7388_22513# m1_7388_22513# m1_6988_22402# m1_7522_21786# m1_7522_21786#
+ pfet$350
Xpfet$348_101 vdd vdd m1_28010_25858# m1_21590_21786# pfet$348
Xnfet$372_16 m1_23486_19550# m1_23486_19550# vss vss m1_23924_20470# vss nfet$372
Xnfet$397_13 fin vss m1_n4623_25487# vss nfet$397
Xnfet$392_6 m1_27190_17836# m1_28113_15778# m1_27292_16202# vss nfet$392
Xnfet$378_4 m1_n789_25858# vss m1_1607_24542# vss nfet$378
Xnfet$373_81 m1_13198_17714# vss m1_10299_17343# vss nfet$373
Xnfet$373_70 m1_n7513_20152# vss m1_18310_16080# vss nfet$373
Xnfet$376_1 sd2 vss m1_21880_15478# vss nfet$376
Xnfet$383_2 m1_17939_22513# m1_17939_22513# vss vss m1_31771_20470# vss nfet$383
Xnfet$390_3 m1_8137_20152# m1_8137_20152# m1_6107_19404# m1_6107_19404# m1_6971_20470#
+ vss nfet$390
Xnfet$369_0 m1_4509_24346# m1_4509_24346# vss vss m1_3991_24542# vss nfet$369
Xnfet$389_25 m1_14743_16202# m1_14743_16202# vss vss m1_14225_16398# vss nfet$389
Xnfet$389_14 m1_n2605_16080# m1_n2605_16080# m1_n3064_17714# m1_n3064_17714# m1_n2507_16398#
+ vss nfet$389
Xpfet$354_8 vdd vdd m1_n1133_19550# m1_n7383_17599# pfet$354
Xnfet$370_82 m1_11415_25662# m1_12259_24224# m1_13363_25658# vss nfet$370
Xnfet$370_71 m1_28147_25662# m1_28371_23922# m1_28635_24542# vss nfet$370
Xnfet$370_60 pd6 vss m1_16322_21786# vss nfet$370
Xpfet$352_12 vdd vdd m1_16452_21590# m1_16322_21786# pfet$352
Xpfet$373_0 vdd vdd m1_n4485_20152# m1_n3822_20130# pfet$373
Xnfet$375_16 m1_17381_17714# vss m1_19969_19550# vss nfet$375
Xnfet$401_0 m1_n8283_20611# vss m1_n8283_19850# vss nfet$401
Xpfet$352_5 vdd vdd m1_1120_21786# m1_488_21786# pfet$352
Xpfet$350_2 vdd m1_7388_22513# m1_7388_22513# m1_6360_22102# m1_8154_21786# m1_8154_21786#
+ pfet$350
Xpfet$348_102 vdd m1_28371_23922# m1_28635_24542# m1_28010_25858# pfet$348
Xpfet$374_10 vdd vdd m1_n10933_25858# fin pfet$374
Xnfet$372_17 m1_12935_19550# m1_12935_19550# vss vss m1_13373_20470# vss nfet$372
Xnfet$399_0 m1_n10933_25858# m1_n8848_25658# m1_n8055_24542# vss nfet$399
Xnfet$392_7 m1_27190_17836# m1_28470_16080# m1_28003_18030# vss nfet$392
Xnfet$378_5 m1_n789_25858# vss m1_488_21786# vss nfet$378
Xnfet$373_82 m1_10299_17343# vss m1_10458_17836# vss nfet$373
Xnfet$373_71 m1_14641_17836# m1_15921_16080# m1_15454_18030# vss nfet$373
Xnfet$373_60 m1_18665_17343# vss m1_18824_17836# vss nfet$373
Xnfet$376_2 sd1 vss m1_26063_15478# vss nfet$376
Xnfet$383_3 m1_24973_22513# m1_24973_22513# vss vss m1_30492_20470# vss nfet$383
Xnfet$390_4 m1_965_15478# m1_965_15478# m1_6107_19404# m1_6107_19404# m1_6339_20470#
+ vss nfet$390
Xnfet$369_1 m1_3893_24224# m1_3893_24224# m1_3537_24542# m1_3537_24542# m1_3991_24542#
+ vss nfet$369
Xnfet$389_26 m1_14127_16080# m1_14127_16080# m1_13668_17714# m1_13668_17714# m1_14225_16398#
+ vss nfet$389
Xpfet$354_9 vdd vdd m1_27003_19550# m1_25747_17714# pfet$354
Xnfet$389_15 m1_n1989_16202# m1_n1989_16202# vss vss m1_n2507_16398# vss nfet$389
Xnfet$381_0 m1_n290_24224# m1_n290_24224# m1_n646_24542# m1_n646_24542# m1_n192_24542#
+ vss nfet$381
Xnfet$370_72 m1_23827_25858# m1_25912_25658# m1_26705_24542# vss nfet$370
Xnfet$370_61 m1_23964_25662# m1_24808_24224# m1_25912_25658# vss nfet$370
Xnfet$370_50 m1_n7513_20152# vss m1_21241_24346# vss nfet$370
Xpfet$352_13 vdd vdd m1_15188_21786# m1_14556_21786# pfet$352
Xpfet$366_0 vdd vdd m1_n7247_17714# m1_n6788_16080# pfet$366
Xpfet$373_1 vdd m1_n4485_21904# vdd m1_9624_19404# pfet$373
Xnfet$375_17 m1_21880_15478# vss m1_25722_20152# vss nfet$375
Xnfet$401_1 m1_n7513_20152# m1_n8283_19850# vss vss nfet$401
Xpfet$352_6 vdd vdd m1_5901_21590# m1_5771_21786# pfet$352
Xpfet$348_103 vdd vdd m1_28635_24542# m1_28991_24224# pfet$348
Xpfet$350_3 vdd m1_9645_21447# m1_9645_21447# m1_10505_22402# m1_11039_21786# m1_11039_21786#
+ pfet$350
Xnfet$399_1 m1_n10796_25662# m1_n10572_23922# m1_n10308_24542# vss nfet$399
Xpfet$374_11 vdd vdd m1_n9336_24346# vss pfet$374
Xnfet$378_6 m1_n910_23922# vss m1_n290_24224# vss nfet$378
Xnfet$373_72 m1_17851_17714# vss m1_18441_17518# vss nfet$373
Xnfet$373_61 m1_20104_16080# vss m1_19747_15778# vss nfet$373
Xnfet$373_50 m1_25747_17714# vss m1_22848_17343# vss nfet$373
Xnfet$383_4 m1_32818_20470# m1_32818_20470# vss vss m1_34329_20470# vss nfet$383
Xnfet$369_2 m1_4997_25658# m1_4997_25658# vss vss m1_5456_25502# vss nfet$369
Xnfet$390_5 m1_5148_15478# m1_5148_15478# m1_9624_19404# m1_9624_19404# m1_9856_20470#
+ vss nfet$390
Xnfet$381_1 m1_814_25658# m1_814_25658# vss vss m1_1273_25502# vss nfet$381
Xnfet$370_73 m1_24309_25858# vss m1_21590_21786# vss nfet$370
Xnfet$370_62 m1_24188_23922# vss m1_24808_24224# vss nfet$370
Xnfet$370_51 m1_19644_25858# m1_21729_25658# m1_22522_24542# vss nfet$370
Xnfet$370_40 m1_15598_25662# m1_16442_24224# m1_17546_25658# vss nfet$370
Xnfet$389_27 m1_18310_16080# m1_18310_16080# vss vss m1_19873_17358# vss nfet$389
Xnfet$389_16 m1_19747_15778# m1_19747_15778# m1_19637_18030# m1_19637_18030# m1_19873_17358#
+ vss nfet$389
Xpfet$359_0 vdd m1_31535_19792# vdd m1_17939_22513# pfet$359
Xpfet$366_1 vdd m1_n7247_17714# vdd m1_n6172_16202# pfet$366
Xnfet$374_0 m1_n1263_21786# vss m1_n1133_21590# vss nfet$374
Xpfet$373_2 vdd m1_n5227_21418# vdd m1_2590_19404# pfet$373
Xpfet$352_14 vdd vdd m1_19969_21590# m1_19839_21786# pfet$352
Xnfet$401_2 m1_n8145_21908# vss m1_n8283_20611# vss nfet$401
Xpfet$352_7 vdd vdd m1_4637_21786# m1_4005_21786# pfet$352
Xpfet$348_104 vdd m1_25912_25658# m1_26705_24542# m1_23964_25662# pfet$348
Xpfet$350_4 vdd vdd vdd m1_9877_22102# m1_9418_21590# m1_9418_21590# pfet$350
Xnfet$399_2 m1_n10933_25858# m1_n10309_25662# m1_n10572_23922# vss nfet$399
Xpfet$374_12 vdd vdd m1_n7082_23622# m1_n8625_26174# pfet$374
Xpfet$348_90 vdd vdd m1_24309_25858# m1_25424_24346# pfet$348
Xnfet$378_7 m1_25107_21786# vss m1_32193_25858# vss nfet$378
Xnfet$373_73 m1_13668_17714# vss m1_16538_15778# vss nfet$373
Xnfet$373_62 m1_18665_17343# m1_20721_15778# m1_20104_16080# vss nfet$373
Xnfet$373_51 m1_n7513_20152# vss m1_22493_16080# vss nfet$373
Xnfet$373_40 m1_n2250_17343# m1_n194_15778# m1_n811_16080# vss nfet$373
Xnfet$383_5 m1_32818_21586# m1_32818_21586# m1_34093_19792# m1_34093_19792# m1_34329_20470#
+ vss nfet$383
Xnfet$369_3 m1_4509_24346# m1_4509_24346# m1_3394_25858# m1_3394_25858# m1_5456_25502#
+ vss nfet$369
Xnfet$390_6 m1_11654_20152# m1_11654_20152# m1_9624_19404# m1_9624_19404# m1_10488_20470#
+ vss nfet$390
Xnfet$370_52 m1_20126_25858# vss m1_22522_24542# vss nfet$370
Xnfet$370_41 pd5 vss m1_12805_21786# vss nfet$370
Xnfet$370_30 m1_n7513_20152# vss m1_17058_24346# vss nfet$370
Xnfet$389_17 m1_22493_16080# m1_22493_16080# vss vss m1_24056_17358# vss nfet$389
Xnfet$381_2 m1_326_24346# m1_326_24346# m1_n789_25858# m1_n789_25858# m1_1273_25502#
+ vss nfet$381
Xpfet$366_2 vdd vdd m1_n5461_18030# m1_n5351_15778# pfet$366
Xpfet$373_3 vdd vdd m1_n5227_21418# m1_6107_19404# pfet$373
Xnfet$374_1 m1_11039_21786# vss m1_11671_21786# vss nfet$374
Xnfet$370_74 pd8 vss m1_23356_21786# vss nfet$370
Xpfet$352_15 vdd vdd m1_27003_21590# m1_26873_21786# pfet$352
Xnfet$370_63 m1_14556_21786# vss m1_19644_25858# vss nfet$370
Xpfet$359_1 vdd vdd m1_30256_19792# m1_21456_22513# pfet$359
Xnfet$401_3 m1_n8283_19850# m1_n8283_20611# vss vss nfet$401
Xpfet$352_8 vdd vdd m1_2384_21590# m1_2254_21786# pfet$352
Xpfet$371_0 vdd vdd m1_n7320_25516# m1_n7186_25858# pfet$371
Xpfet$348_105 vdd vdd m1_30888_24542# m1_28492_25858# pfet$348
Xpfet$350_5 vdd m1_9645_21447# m1_9645_21447# m1_9877_22102# m1_11671_21786# m1_11671_21786#
+ pfet$350
Xpfet$374_13 vdd vdd m1_n8055_24542# m1_n8625_26174# pfet$374
Xpfet$348_91 vdd vdd m1_23356_21786# pd8 pfet$348
Xpfet$348_80 vdd vdd m1_17058_24346# m1_n7513_20152# pfet$348
Xnfet$399_3 m1_n10796_25662# m1_n9952_24224# m1_n8848_25658# vss nfet$399
Xnfet$378_8 m1_32193_25858# vss m1_32330_25662# vss nfet$378
Xnfet$397_0 m1_n8625_26174# vss m1_n8055_24542# vss nfet$397
Xnfet$373_74 m1_14482_17343# vss m1_14641_17836# vss nfet$373
Xnfet$373_63 m1_13668_17714# vss m1_14258_17518# vss nfet$373
Xnfet$373_52 m1_23007_17836# m1_24287_16080# m1_23820_18030# vss nfet$373
Xnfet$373_30 sd6 vss m1_5148_15478# vss nfet$373
Xnfet$373_41 m1_n2091_17836# m1_n1168_15778# m1_n1989_16202# vss nfet$373
Xnfet$383_6 m1_354_22513# m1_354_22513# m1_31535_22102# m1_31535_22102# m1_31771_21430#
+ vss nfet$383
Xnfet$390_7 m1_n7401_15478# m1_n7401_15478# m1_n927_19404# m1_n927_19404# m1_n695_20470#
+ vss nfet$390
Xnfet$369_4 m1_12259_24224# m1_12259_24224# m1_11903_24542# m1_11903_24542# m1_12357_24542#
+ vss nfet$369
Xnfet$389_18 m1_23930_15778# m1_23930_15778# m1_23820_18030# m1_23820_18030# m1_24056_17358#
+ vss nfet$389
Xnfet$381_3 m1_326_24346# m1_326_24346# vss vss m1_n192_24542# vss nfet$381
Xnfet$374_2 m1_12805_21786# vss m1_12935_21590# vss nfet$374
Xnfet$370_75 m1_28371_23922# vss m1_28991_24224# vss nfet$370
Xpfet$352_16 vdd vdd m1_29256_21786# m1_28624_21786# pfet$352
Xnfet$370_64 m1_19644_25858# vss m1_19781_25662# vss nfet$370
Xnfet$370_53 m1_23827_25858# m1_24451_25662# m1_24188_23922# vss nfet$370
Xnfet$370_42 m1_15943_25858# vss m1_16085_25662# vss nfet$370
Xnfet$370_31 m1_15943_25858# vss m1_18339_24542# vss nfet$370
Xpfet$359_2 vdd m1_30256_19792# vdd m1_24973_22513# pfet$359
Xnfet$370_20 pd3 vss m1_5771_21786# vss nfet$370
Xpfet$366_3 vdd m1_n5461_18030# vdd m1_n6788_16080# pfet$366
Xpfet$373_4 vdd vdd m1_n4485_21904# m1_n3822_21786# pfet$373
Xpfet$364_0 vdd vdd fout m1_34093_22102# pfet$364
Xpfet$352_9 vdd vdd m1_22222_21786# m1_21590_21786# pfet$352
Xpfet$371_1 vdd vdd m1_n6111_25858# m1_n6856_24542# pfet$371
Xpfet$350_6 vdd vdd vdd m1_10505_22402# m1_9288_21786# m1_9288_21786# pfet$350
Xpfet$348_106 vdd vdd m1_25107_21786# m1_28492_25858# pfet$348
Xpfet$348_92 vdd vdd m1_28492_25858# m1_29607_24346# pfet$348
Xpfet$348_81 vdd vdd m1_18339_24542# m1_15943_25858# pfet$348
Xpfet$348_70 vdd vdd m1_14156_24542# m1_11760_25858# pfet$348
Xnfet$399_4 m1_n4623_25487# m1_n2567_23922# m1_n3184_24224# vss nfet$399
Xnfet$378_9 m1_n7513_20152# vss m1_33790_24346# vss nfet$378
Xnfet$373_75 sd3 vss m1_17697_15478# vss nfet$373
Xnfet$373_64 m1_13668_17714# vss m1_13198_17714# vss nfet$373
Xnfet$373_53 m1_22848_17343# vss m1_23007_17836# vss nfet$373
Xnfet$373_31 m1_1933_17343# m1_3989_15778# m1_3372_16080# vss nfet$373
Xnfet$373_20 m1_1119_17714# vss m1_1709_17518# vss nfet$373
Xnfet$373_42 m1_n811_16080# vss m1_n1168_15778# vss nfet$373
Xnfet$397_1 m1_n8625_26174# vss m1_n7082_23622# vss nfet$397
Xnfet$383_7 m1_3871_22513# m1_3871_22513# vss vss m1_31771_21430# vss nfet$383
Xnfet$390_8 m1_26063_15478# m1_26063_15478# m1_n3822_20130# m1_n3822_20130# m1_27441_20470#
+ vss nfet$390
Xnfet$369_5 m1_8692_24346# m1_8692_24346# vss vss m1_8174_24542# vss nfet$369
Xnfet$381_4 m1_33174_24224# m1_33174_24224# m1_32818_24542# m1_32818_24542# m1_33272_24542#
+ vss nfet$381
Xnfet$389_19 m1_23109_16202# m1_23109_16202# vss vss m1_22591_16398# vss nfet$389
Xnfet$374_3 m1_9288_21786# vss m1_9418_21590# vss nfet$374
Xpfet$352_17 vdd vdd m1_25739_21786# m1_25107_21786# pfet$352
Xnfet$370_76 m1_28492_25858# vss m1_28634_25662# vss nfet$370
Xnfet$370_65 m1_28492_25858# vss m1_25107_21786# vss nfet$370
Xnfet$370_54 m1_24309_25858# vss m1_24451_25662# vss nfet$370
Xnfet$370_43 m1_15461_25858# vss m1_15598_25662# vss nfet$370
Xnfet$370_32 m1_15461_25858# m1_17546_25658# m1_18339_24542# vss nfet$370
Xpfet$359_3 vdd vdd m1_34843_21786# m1_34093_19792# pfet$359
Xpfet$366_4 vdd vdd m1_26217_17714# m1_26676_16080# pfet$366
Xnfet$370_21 m1_11278_25858# m1_11902_25662# m1_11639_23922# vss nfet$370
Xnfet$370_10 m1_7577_25858# vss m1_9973_24542# vss nfet$370
Xpfet$373_5 vdd m1_n6839_21786# vdd m1_n5764_21786# pfet$373
Xnfet$372_0 m1_n3534_17714# m1_n3534_17714# vss vss m1_3454_20470# vss nfet$372
Xpfet$357_0 vdd vdd m1_n646_24542# m1_n290_24224# pfet$357
Xpfet$350_7 vdd m1_354_22513# m1_354_22513# m1_n674_22102# m1_1120_21786# m1_1120_21786#
+ pfet$350
Xpfet$348_107 vdd m1_24309_25858# vdd m1_25912_25658# pfet$348
Xpfet$348_93 vdd m1_28991_24224# m1_30095_25658# m1_28010_25858# pfet$348
Xpfet$348_82 vdd vdd m1_21241_24346# m1_n7513_20152# pfet$348
Xpfet$348_71 vdd vdd m1_11039_21786# m1_11760_25858# pfet$348
Xpfet$348_60 vdd vdd m1_20126_25858# m1_21241_24346# pfet$348
Xnfet$399_5 m1_n4464_25980# m1_n3541_23922# m1_n4362_24346# vss nfet$399
Xnfet$373_76 m1_14482_17343# m1_16538_15778# m1_15921_16080# vss nfet$373
Xnfet$373_65 m1_14482_17343# m1_14743_16202# m1_14258_17518# vss nfet$373
Xnfet$373_54 m1_22848_17343# m1_23109_16202# m1_22624_17518# vss nfet$373
Xnfet$373_32 m1_2092_17836# m1_3015_15778# m1_2194_16202# vss nfet$373
Xnfet$373_21 m1_1933_17343# m1_2194_16202# m1_1709_17518# vss nfet$373
Xnfet$373_10 m1_11738_16080# vss m1_11381_15778# vss nfet$373
Xnfet$373_43 sd8 vss m1_n3218_15478# vss nfet$373
Xnfet$397_2 vss vss m1_n9336_24346# vss nfet$397
Xnfet$390_9 m1_29239_20152# m1_29239_20152# m1_n3822_20130# m1_n3822_20130# m1_28073_20470#
+ vss nfet$390
Xnfet$369_6 m1_8076_24224# m1_8076_24224# m1_7720_24542# m1_7720_24542# m1_8174_24542#
+ vss nfet$369
Xnfet$381_5 m1_33790_24346# m1_33790_24346# vss vss m1_33272_24542# vss nfet$381
Xnfet$374_4 m1_7522_21786# vss m1_8154_21786# vss nfet$374
Xnfet$370_77 m1_28010_25858# vss m1_28147_25662# vss nfet$370
Xnfet$370_66 m1_28010_25858# m1_30095_25658# m1_30888_24542# vss nfet$370
Xnfet$370_55 m1_23827_25858# vss m1_23964_25662# vss nfet$370
Xnfet$370_44 m1_15822_23922# vss m1_16442_24224# vss nfet$370
Xnfet$370_33 m1_11760_25858# vss m1_14156_24542# vss nfet$370
Xpfet$359_4 vdd m1_34093_19792# vdd m1_32818_20470# pfet$359
Xpfet$366_5 vdd m1_26217_17714# vdd m1_27292_16202# pfet$366
Xnfet$370_22 m1_11760_25858# vss m1_11902_25662# vss nfet$370
Xnfet$370_11 m1_7522_21786# vss m1_11278_25858# vss nfet$370
Xpfet$373_6 vdd vdd m1_n6973_21481# m1_n6839_21786# pfet$373
Xnfet$372_1 m1_2384_19550# m1_2384_19550# vss vss m1_2822_20470# vss nfet$372
Xpfet$357_1 vdd m1_n789_25858# vdd m1_814_25658# pfet$357
Xpfet$348_108 vdd vdd m1_25424_24346# m1_n7513_20152# pfet$348
Xpfet$350_8 vdd vdd vdd m1_6360_22102# m1_5901_21590# m1_5901_21590# pfet$350
Xpfet$348_94 vdd m1_28492_25858# vdd m1_30095_25658# pfet$348
Xpfet$348_83 vdd m1_21729_25658# m1_22522_24542# m1_19781_25662# pfet$348
Xpfet$348_72 vdd m1_13363_25658# m1_14156_24542# m1_11415_25662# pfet$348
Xpfet$348_61 vdd m1_24452_24542# vdd m1_25424_24346# pfet$348
Xpfet$348_50 vdd vdd m1_20268_25662# m1_20126_25858# pfet$348
Xnfet$399_6 m1_n4464_25980# m1_n3184_24224# m1_n3651_26174# vss nfet$399
Xnfet$397_3 fin vss m1_n10933_25858# vss nfet$397
Xnfet$373_77 sd4 vss m1_13514_15478# vss nfet$373
Xnfet$373_66 m1_n7513_20152# vss m1_14127_16080# vss nfet$373
Xnfet$373_55 m1_22034_17714# vss m1_24904_15778# vss nfet$373
Xnfet$373_44 m1_n2091_17836# m1_n811_16080# m1_n1278_18030# vss nfet$373
Xnfet$373_33 sd7 vss m1_965_15478# vss nfet$373
Xnfet$373_22 m1_6116_17343# m1_6377_16202# m1_5892_17518# vss nfet$373
Xnfet$373_11 m1_10299_17343# m1_12355_15778# m1_11738_16080# vss nfet$373
Xnfet$369_7 m1_9180_25658# m1_9180_25658# vss vss m1_9639_25502# vss nfet$369
Xnfet$395_0 m1_n7082_23622# m1_n6856_24542# vss vss nfet$395
Xnfet$381_6 m1_33790_24346# m1_33790_24346# m1_32675_25947# m1_32675_25947# m1_34737_25502#
+ vss nfet$381
Xnfet$370_78 m1_28010_25858# m1_28634_25662# m1_28371_23922# vss nfet$370
Xnfet$370_67 m1_28492_25858# vss m1_30888_24542# vss nfet$370
Xnfet$370_56 m1_19781_25662# m1_20625_24224# m1_21729_25658# vss nfet$370
Xnfet$370_45 m1_15461_25858# m1_16085_25662# m1_15822_23922# vss nfet$370
Xnfet$370_34 m1_11278_25858# m1_13363_25658# m1_14156_24542# vss nfet$370
Xpfet$366_6 vdd vdd m1_28003_18030# m1_28113_15778# pfet$366
Xpfet$359_5 vdd vdd m1_34093_19792# m1_32818_21586# pfet$359
Xnfet$370_23 m1_11278_25858# vss m1_11415_25662# vss nfet$370
Xnfet$370_12 m1_7577_25858# vss m1_7522_21786# vss nfet$370
Xpfet$373_7 vdd vdd m1_n6839_21786# m1_n6380_21786# pfet$373
Xnfet$374_5 m1_488_21786# vss m1_1120_21786# vss nfet$374
Xnfet$372_2 m1_5901_19550# m1_5901_19550# vss vss m1_6339_20470# vss nfet$372
Xpfet$357_2 vdd vdd m1_n789_25858# m1_326_24346# pfet$357
Xpfet$348_109 vdd m1_12259_24224# m1_13363_25658# m1_11278_25858# pfet$348
Xpfet$350_9 vdd m1_3871_22513# m1_3871_22513# m1_3471_22402# m1_4005_21786# m1_4005_21786#
+ pfet$350
Xpfet$362_0 vdd m1_34093_22102# vdd m1_28490_22513# pfet$362
Xnfet$399_7 m1_n4623_25487# m1_n4362_24346# m1_n4847_25662# vss nfet$399
Xpfet$348_95 vdd vdd m1_28991_24224# m1_28371_23922# pfet$348
Xpfet$348_84 vdd vdd m1_23827_25858# m1_18073_21786# pfet$348
Xpfet$348_73 vdd m1_16086_24542# vdd m1_17058_24346# pfet$348
Xpfet$348_62 vdd vdd m1_24452_24542# m1_24808_24224# pfet$348
Xpfet$348_51 vdd vdd m1_20625_24224# m1_20005_23922# pfet$348
Xpfet$348_40 vdd vdd m1_11760_25858# m1_12875_24346# pfet$348
Xpfet$350_30 vdd vdd vdd m1_17539_22402# m1_16322_21786# m1_16322_21786# pfet$350
Xnfet$397_4 m1_n10572_23922# vss m1_n9952_24224# vss nfet$397
Xnfet$373_78 m1_14641_17836# m1_15564_15778# m1_14743_16202# vss nfet$373
Xnfet$373_67 m1_17381_17714# vss m1_14482_17343# vss nfet$373
Xnfet$373_56 m1_24287_16080# vss m1_23930_15778# vss nfet$373
Xnfet$373_45 m1_n3064_17714# vss m1_n194_15778# vss nfet$373
Xnfet$373_34 m1_n2250_17343# vss m1_n2091_17836# vss nfet$373
Xnfet$373_23 m1_5302_17714# vss m1_4832_17714# vss nfet$373
Xnfet$373_12 m1_9485_17714# vss m1_12355_15778# vss nfet$373
Xnfet$369_8 m1_8692_24346# m1_8692_24346# m1_7577_25858# m1_7577_25858# m1_9639_25502#
+ vss nfet$369
Xnfet$388_0 fout vss m1_35837_22102# vss nfet$388
Xnfet$395_1 m1_n8283_19850# vss m1_n6856_24542# vss nfet$395
Xnfet$381_7 m1_34278_25658# m1_34278_25658# vss vss m1_34737_25502# vss nfet$381
Xnfet$370_57 m1_20126_25858# vss m1_20268_25662# vss nfet$370
Xnfet$370_46 m1_20126_25858# vss m1_18073_21786# vss nfet$370
Xnfet$370_35 m1_15598_25662# m1_15822_23922# m1_16086_24542# vss nfet$370
Xpfet$366_7 vdd m1_28003_18030# vdd m1_26676_16080# pfet$366
Xnfet$370_24 m1_7095_25858# m1_7719_25662# m1_7456_23922# vss nfet$370
Xnfet$370_13 m1_11415_25662# m1_11639_23922# m1_11903_24542# vss nfet$370
Xnfet$374_6 m1_5771_21786# vss m1_5901_21590# vss nfet$374
Xnfet$370_79 pd7 vss m1_19839_21786# vss nfet$370
Xnfet$370_68 m1_n7513_20152# vss m1_29607_24346# vss nfet$370
Xpfet$359_6 vdd vdd m1_31535_19792# m1_14422_22513# pfet$359
Xnfet$372_3 m1_4832_17714# m1_4832_17714# vss vss m1_10488_20470# vss nfet$372
Xpfet$357_3 vdd m1_n646_24542# vdd m1_326_24346# pfet$357
Xnfet$370_0 m1_3394_25858# vss m1_5790_24542# vss nfet$370
Xpfet$362_1 vdd vdd m1_34093_22102# m1_34843_21786# pfet$362
Xpfet$355_0 vdd vdd m1_n7401_15478# sd9 pfet$355
Xpfet$348_96 vdd m1_28635_24542# vdd m1_29607_24346# pfet$348
Xpfet$348_85 vdd m1_24188_23922# m1_24452_24542# m1_23827_25858# pfet$348
Xpfet$348_74 vdd vdd m1_14556_21786# m1_15943_25858# pfet$348
Xpfet$348_63 vdd vdd m1_19781_25662# m1_19644_25858# pfet$348
Xpfet$348_52 vdd m1_20268_25662# m1_20005_23922# m1_19781_25662# pfet$348
Xpfet$348_41 vdd vdd m1_9288_21786# pd4 pfet$348
Xpfet$348_30 vdd vdd m1_2912_25858# m1_488_21786# pfet$348
Xpfet$350_31 vdd vdd vdd m1_27462_22102# m1_27003_21590# m1_27003_21590# pfet$350
Xpfet$350_20 vdd vdd vdd m1_20428_22102# m1_19969_21590# m1_19969_21590# pfet$350
Xnfet$397_5 m1_n10933_25858# vss m1_n10796_25662# vss nfet$397
Xnfet$373_79 m1_15921_16080# vss m1_15564_15778# vss nfet$373
Xnfet$373_68 m1_18665_17343# m1_18926_16202# m1_18441_17518# vss nfet$373
Xnfet$373_57 m1_22848_17343# m1_24904_15778# m1_24287_16080# vss nfet$373
Xnfet$373_46 m1_22034_17714# vss m1_21564_17714# vss nfet$373
Xnfet$373_24 m1_4832_17714# vss m1_1933_17343# vss nfet$373
Xnfet$373_13 m1_10458_17836# m1_11381_15778# m1_10560_16202# vss nfet$373
Xnfet$373_35 m1_n7513_20152# vss m1_5761_16080# vss nfet$373
Xnfet$369_9 m1_17058_24346# m1_17058_24346# vss vss m1_16540_24542# vss nfet$369
Xnfet$388_1 define m1_35837_22102# vss vss nfet$388
Xnfet$374_7 m1_4005_21786# vss m1_4637_21786# vss nfet$374
Xpfet$359_7 vdd vdd m1_31535_22102# m1_354_22513# pfet$359
Xnfet$370_69 m1_24309_25858# vss m1_26705_24542# vss nfet$370
Xnfet$370_58 m1_20005_23922# vss m1_20625_24224# vss nfet$370
Xnfet$370_47 m1_23964_25662# m1_24188_23922# m1_24452_24542# vss nfet$370
Xnfet$370_36 m1_11760_25858# vss m1_11039_21786# vss nfet$370
Xnfet$370_25 m1_7232_25662# m1_8076_24224# m1_9180_25658# vss nfet$370
Xnfet$370_14 m1_n7513_20152# vss m1_8692_24346# vss nfet$370
Xpfet$357_4 vdd vdd m1_32675_25947# m1_33790_24346# pfet$357
Xnfet$372_4 m1_9418_19550# m1_9418_19550# vss vss m1_9856_20470# vss nfet$372
Xnfet$370_1 m1_2912_25858# m1_4997_25658# m1_5790_24542# vss nfet$370
Xpfet$362_2 vdd vdd m1_30256_22102# m1_7388_22513# pfet$362
Xpfet$355_1 vdd vdd m1_21880_15478# sd2 pfet$355
Xpfet$348_0 vdd vdd m1_3049_25662# m1_2912_25858# pfet$348
Xpfet$348_97 vdd vdd m1_21590_21786# m1_24309_25858# pfet$348
Xpfet$348_86 vdd m1_28634_25662# m1_28371_23922# m1_28147_25662# pfet$348
Xpfet$348_75 vdd vdd m1_19644_25858# m1_14556_21786# pfet$348
Xpfet$348_64 vdd vdd m1_22522_24542# m1_20126_25858# pfet$348
Xpfet$348_53 vdd m1_20625_24224# m1_21729_25658# m1_19644_25858# pfet$348
Xpfet$348_42 vdd m1_11760_25858# vdd m1_13363_25658# pfet$348
Xpfet$348_31 vdd m1_3273_23922# m1_3537_24542# m1_2912_25858# pfet$348
Xpfet$348_20 vdd vdd m1_4509_24346# m1_n7513_20152# pfet$348
Xpfet$350_32 vdd m1_28490_22513# m1_28490_22513# m1_28090_22402# m1_28624_21786# m1_28624_21786#
+ pfet$350
Xpfet$350_21 vdd vdd vdd m1_21056_22402# m1_19839_21786# m1_19839_21786# pfet$350
Xpfet$350_10 vdd m1_3871_22513# m1_3871_22513# m1_2843_22102# m1_4637_21786# m1_4637_21786#
+ pfet$350
Xnfet$373_69 m1_17851_17714# vss m1_17381_17714# vss nfet$373
Xnfet$373_58 m1_23007_17836# m1_23930_15778# m1_23109_16202# vss nfet$373
Xnfet$373_47 m1_22034_17714# vss m1_22624_17518# vss nfet$373
Xnfet$373_25 m1_2092_17836# m1_3372_16080# m1_2905_18030# vss nfet$373
Xnfet$373_14 m1_6116_17343# m1_8172_15778# m1_7555_16080# vss nfet$373
Xnfet$373_36 m1_n3064_17714# vss m1_n2474_17518# vss nfet$373
Xnfet$397_6 m1_n10452_25858# vss m1_n10309_25662# vss nfet$397
Xnfet$374_8 m1_2254_21786# vss m1_2384_21590# vss nfet$374
Xnfet$370_59 m1_19644_25858# m1_20268_25662# m1_20005_23922# vss nfet$370
Xnfet$370_48 m1_18073_21786# vss m1_23827_25858# vss nfet$370
Xnfet$370_37 m1_11039_21786# vss m1_15461_25858# vss nfet$370
Xnfet$370_26 m1_7095_25858# m1_9180_25658# m1_9973_24542# vss nfet$370
Xnfet$370_15 m1_7232_25662# m1_7456_23922# m1_7720_24542# vss nfet$370
Xnfet$393_0 m1_n5351_15778# m1_n5351_15778# m1_n5461_18030# m1_n5461_18030# m1_n5225_17358#
+ vss nfet$393
Xpfet$378_0 vdd vdd m1_n5227_20152# m1_n2543_20130# pfet$378
Xnfet$372_5 m1_649_17714# m1_649_17714# vss vss m1_6971_20470# vss nfet$372
Xpfet$357_5 vdd m1_32675_25947# vdd m1_34278_25658# pfet$357
Xpfet$353_10 vdd vdd m1_27031_17343# m1_n10452_25858# pfet$353
Xnfet$370_2 m1_n7513_20152# vss m1_4509_24346# vss nfet$370
Xpfet$355_2 vdd vdd m1_26063_15478# sd1 pfet$355
Xpfet$362_3 vdd m1_31535_22102# vdd m1_3871_22513# pfet$362
Xpfet$348_1 vdd m1_3536_25662# m1_3273_23922# m1_3049_25662# pfet$348
Xpfet$348_98 vdd m1_30095_25658# m1_30888_24542# m1_28147_25662# pfet$348
Xpfet$348_87 vdd vdd m1_28147_25662# m1_28010_25858# pfet$348
Xpfet$348_76 vdd m1_20005_23922# m1_20269_24542# m1_19644_25858# pfet$348
Xpfet$348_65 vdd vdd m1_18073_21786# m1_20126_25858# pfet$348
Xpfet$348_54 vdd vdd m1_24808_24224# m1_24188_23922# pfet$348
Xpfet$348_43 vdd vdd m1_12805_21786# pd5 pfet$348
Xpfet$348_32 vdd vdd m1_7720_24542# m1_8076_24224# pfet$348
Xpfet$348_21 vdd m1_7456_23922# m1_7720_24542# m1_7095_25858# pfet$348
Xpfet$348_10 vdd m1_8076_24224# m1_9180_25658# m1_7095_25858# pfet$348
Xpfet$350_33 vdd m1_28490_22513# m1_28490_22513# m1_27462_22102# m1_29256_21786# m1_29256_21786#
+ pfet$350
Xpfet$350_22 vdd m1_21456_22513# m1_21456_22513# m1_20428_22102# m1_22222_21786# m1_22222_21786#
+ pfet$350
Xpfet$360_0 vdd m1_n647_25662# m1_n910_23922# m1_n1134_25662# pfet$360
Xpfet$350_11 vdd vdd vdd m1_2843_22102# m1_2384_21590# m1_2384_21590# pfet$350
Xnfet$373_59 m1_17851_17714# vss m1_20721_15778# vss nfet$373
Xnfet$373_48 m1_18824_17836# m1_20104_16080# m1_19637_18030# vss nfet$373
Xnfet$373_26 m1_5302_17714# vss m1_5892_17518# vss nfet$373
Xnfet$373_15 m1_5302_17714# vss m1_8172_15778# vss nfet$373
Xnfet$373_37 m1_n7513_20152# vss m1_n2605_16080# vss nfet$373
Xnfet$397_7 m1_n7320_25516# vss m1_n2567_23922# vss nfet$397
Xpfet$356_10 vdd vdd m1_35071_24542# m1_32675_25947# pfet$356
Xnfet$374_9 m1_23356_21786# vss m1_23486_21590# vss nfet$374
Xnfet$370_49 m1_19781_25662# m1_20005_23922# m1_20269_24542# vss nfet$370
Xnfet$370_38 m1_n7513_20152# vss m1_12875_24346# vss nfet$370
Xnfet$386_0 m1_34093_19792# vss m1_34843_21786# vss nfet$386
Xnfet$370_27 m1_7577_25858# vss m1_7719_25662# vss nfet$370
Xnfet$370_16 m1_4005_21786# vss m1_7095_25858# vss nfet$370
Xnfet$393_1 m1_n6788_16080# m1_n6788_16080# vss vss m1_n5225_17358# vss nfet$393
Xpfet$378_1 vdd m1_n4485_20152# vdd m1_n3206_20274# pfet$378
Xnfet$372_6 m1_n1133_19550# m1_n1133_19550# vss vss m1_n695_20470# vss nfet$372
Xpfet$357_6 vdd vdd m1_32818_24542# m1_33174_24224# pfet$357
Xpfet$353_11 vdd vdd m1_26807_17518# m1_26217_17714# pfet$353
Xpfet$362_4 vdd m1_30256_22102# vdd m1_9645_21447# pfet$362
Xnfet$370_3 m1_488_21786# vss m1_2912_25858# vss nfet$370
Xpfet$348_99 vdd vdd m1_26705_24542# m1_24309_25858# pfet$348
Xpfet$348_88 vdd vdd m1_28634_25662# m1_28492_25858# pfet$348
Xpfet$348_77 vdd vdd m1_20269_24542# m1_20625_24224# pfet$348
Xpfet$348_66 vdd vdd m1_15461_25858# m1_11039_21786# pfet$348
Xpfet$348_55 vdd m1_24451_25662# m1_24188_23922# m1_23964_25662# pfet$348
Xpfet$348_44 vdd m1_15943_25858# vdd m1_17546_25658# pfet$348
Xpfet$348_33 vdd vdd m1_7522_21786# m1_7577_25858# pfet$348
Xpfet$348_22 vdd vdd m1_3537_24542# m1_3893_24224# pfet$348
Xpfet$348_11 vdd vdd m1_7719_25662# m1_7577_25858# pfet$348
Xpfet$348_2 vdd vdd m1_3394_25858# m1_4509_24346# pfet$348
Xpfet$353_0 vdd vdd m1_n6274_17836# m1_n6433_17343# pfet$353
Xpfet$360_1 vdd m1_n910_23922# m1_n646_24542# m1_n1271_25858# pfet$360
Xpfet$350_34 vdd vdd vdd m1_28090_22402# m1_26873_21786# m1_26873_21786# pfet$350
Xpfet$350_23 vdd vdd vdd m1_23945_22102# m1_23486_21590# m1_23486_21590# pfet$350
Xnfet$397_8 m1_n4623_25487# vss m1_n4464_25980# vss nfet$397
Xpfet$350_12 vdd vdd vdd m1_3471_22402# m1_2254_21786# m1_2254_21786# pfet$350
Xnfet$373_49 m1_21564_17714# vss m1_18665_17343# vss nfet$373
Xnfet$373_27 m1_1119_17714# vss m1_3989_15778# vss nfet$373
Xnfet$373_16 m1_6275_17836# m1_7198_15778# m1_6377_16202# vss nfet$373
Xnfet$373_38 m1_n2250_17343# m1_n1989_16202# m1_n2474_17518# vss nfet$373
Xpfet$356_11 vdd vdd m1_32817_25662# m1_32675_25947# pfet$356
Xnfet$370_39 pd4 vss m1_9288_21786# vss nfet$370
Xnfet$386_1 m1_30256_19792# vss m1_32818_20470# vss nfet$386
Xnfet$370_28 m1_3394_25858# vss m1_4005_21786# vss nfet$370
Xnfet$370_17 m1_11639_23922# vss m1_12259_24224# vss nfet$370
Xnfet$393_2 m1_n6788_16080# m1_n6788_16080# m1_n7247_17714# m1_n7247_17714# m1_n6690_16398#
+ vss nfet$393
Xnfet$379_0 m1_n1134_25662# m1_n910_23922# m1_n646_24542# vss nfet$379
Xpfet$378_2 vdd m1_n5227_20152# vdd m1_n1927_20274# pfet$378
Xnfet$372_7 m1_n7383_17599# m1_n7383_17599# vss vss m1_n63_20470# vss nfet$372
Xpfet$357_7 vdd m1_32818_24542# vdd m1_33790_24346# pfet$357
Xpfet$353_12 vdd vdd m1_26676_16080# m1_n7513_20152# pfet$353
Xnfet$370_4 m1_2912_25858# vss m1_3049_25662# vss nfet$370
Xpfet$348_34 vdd m1_9180_25658# m1_9973_24542# m1_7232_25662# pfet$348
Xpfet$348_23 vdd m1_3537_24542# vdd m1_4509_24346# pfet$348
Xpfet$348_12 vdd m1_7577_25858# vdd m1_9180_25658# pfet$348
Xpfet$348_3 vdd m1_3394_25858# vdd m1_4997_25658# pfet$348
Xpfet$348_89 vdd vdd m1_19839_21786# pd7 pfet$348
Xpfet$348_78 vdd m1_20269_24542# vdd m1_21241_24346# pfet$348
Xpfet$348_67 vdd m1_15822_23922# m1_16086_24542# m1_15461_25858# pfet$348
Xpfet$348_56 vdd m1_24808_24224# m1_25912_25658# m1_23827_25858# pfet$348
Xpfet$348_45 vdd vdd m1_16442_24224# m1_15822_23922# pfet$348
Xpfet$353_1 vdd vdd m1_n4377_15778# m1_n7247_17714# pfet$353
Xpfet$360_2 vdd m1_n290_24224# m1_814_25658# m1_n1271_25858# pfet$360
Xpfet$350_35 vdd vdd vdd m1_13394_22102# m1_12935_21590# m1_12935_21590# pfet$350
Xpfet$350_24 vdd m1_17939_22513# m1_17939_22513# m1_16911_22102# m1_18705_21786# m1_18705_21786#
+ pfet$350
Xpfet$350_13 vdd vdd vdd m1_6988_22402# m1_5771_21786# m1_5771_21786# pfet$350
Xnfet$397_9 m1_n3184_24224# vss m1_n3541_23922# vss nfet$397
Xnfet$373_28 m1_1933_17343# vss m1_2092_17836# vss nfet$373
Xnfet$373_17 m1_649_17714# vss m1_n2250_17343# vss nfet$373
Xnfet$373_39 m1_n3064_17714# vss m1_n3534_17714# vss nfet$373
Xpfet$356_12 vdd vdd m1_32193_25858# m1_25107_21786# pfet$356
Xnfet$370_29 m1_15943_25858# vss m1_14556_21786# vss nfet$370
Xnfet$370_18 m1_7095_25858# vss m1_7232_25662# vss nfet$370
Xnfet$393_3 m1_n6172_16202# m1_n6172_16202# vss vss m1_n6690_16398# vss nfet$393
Xnfet$386_2 m1_31535_19792# m1_32818_20470# vss vss nfet$386
Xpfet$378_3 vdd m1_n6839_20152# vdd m1_n927_19404# pfet$378
Xnfet$379_1 m1_n1271_25858# m1_n647_25662# m1_n910_23922# vss nfet$379
Xnfet$372_8 m1_27003_19550# m1_27003_19550# vss vss m1_27441_20470# vss nfet$372
Xnfet$391_0 m1_35837_22102# vss m1_n7513_20152# vss nfet$391
Xpfet$353_13 vdd vdd m1_25747_17714# m1_26217_17714# pfet$353
Xpfet$376_0 vdd vdd vdd m1_n8047_19550# m1_n7513_20152# m1_n7513_20152# pfet$376
Xnfet$370_5 m1_2912_25858# m1_3536_25662# m1_3273_23922# vss nfet$370
Xpfet$348_4 vdd vdd m1_3893_24224# m1_3273_23922# pfet$348
Xnfet$404_0 m1_n4485_20152# m1_n6380_21786# vss vss nfet$404
Xpfet$348_79 vdd m1_17546_25658# m1_18339_24542# m1_15598_25662# pfet$348
Xpfet$348_68 vdd vdd m1_16086_24542# m1_16442_24224# pfet$348
Xpfet$348_57 vdd vdd m1_24451_25662# m1_24309_25858# pfet$348
Xpfet$348_46 vdd m1_16442_24224# m1_17546_25658# m1_15461_25858# pfet$348
Xpfet$348_35 vdd m1_7720_24542# vdd m1_8692_24346# pfet$348
Xpfet$348_24 vdd vdd m1_5790_24542# m1_3394_25858# pfet$348
Xpfet$348_13 vdd vdd m1_12259_24224# m1_11639_23922# pfet$348
Xpfet$360_3 vdd m1_814_25658# m1_1607_24542# m1_n1134_25662# pfet$360
Xpfet$353_2 vdd vdd m1_n5351_15778# m1_n4994_16080# pfet$353
Xpfet$350_25 vdd m1_17939_22513# m1_17939_22513# m1_17539_22402# m1_18073_21786# m1_18073_21786#
+ pfet$350
Xpfet$350_14 vdd vdd vdd m1_n46_22402# m1_n1263_21786# m1_n1263_21786# pfet$350
Xnfet$373_29 m1_3372_16080# vss m1_3015_15778# vss nfet$373
Xnfet$373_18 m1_1119_17714# vss m1_649_17714# vss nfet$373
Xpfet$356_13 vdd vdd m1_33790_24346# m1_n7513_20152# pfet$356
Xnfet$386_3 m1_30256_22102# vss m1_32818_21586# vss nfet$386
Xnfet$393_4 m1_28113_15778# m1_28113_15778# m1_28003_18030# m1_28003_18030# m1_28239_17358#
+ vss nfet$393
Xnfet$370_19 m1_7456_23922# vss m1_8076_24224# vss nfet$370
Xpfet$378_4 vdd vdd m1_n6839_20152# m1_n6973_21481# pfet$378
Xnfet$379_2 m1_n1271_25858# m1_814_25658# m1_1607_24542# vss nfet$379
Xnfet$384_0 m1_34843_21786# m1_34843_21786# m1_34093_22102# m1_34093_22102# m1_34329_21430#
+ vss nfet$384
Xnfet$372_9 m1_25747_17714# m1_25747_17714# vss vss m1_28073_20470# vss nfet$372
Xpfet$376_1 vdd m1_n8283_19850# m1_n8283_19850# m1_n8047_19550# m1_n8283_20611# m1_n8283_20611#
+ pfet$376
Xpfet$369_0 vdd vdd vdd m1_n6624_23622# m1_n7082_23622# m1_n7082_23622# pfet$369
Xnfet$370_6 m1_3049_25662# m1_3893_24224# m1_4997_25658# vss nfet$370
Xpfet$348_5 vdd m1_3893_24224# m1_4997_25658# m1_2912_25858# pfet$348
Xnfet$404_1 m1_n5227_20152# vss m1_n6380_21786# vss nfet$404
Xpfet$348_69 vdd vdd m1_12875_24346# m1_n7513_20152# pfet$348
Xpfet$348_58 vdd vdd m1_23964_25662# m1_23827_25858# pfet$348
Xpfet$348_47 vdd vdd m1_15943_25858# m1_17058_24346# pfet$348
Xpfet$348_36 vdd vdd m1_8692_24346# m1_n7513_20152# pfet$348
Xpfet$348_25 vdd vdd m1_4005_21786# m1_3394_25858# pfet$348
Xpfet$348_14 vdd vdd m1_11902_25662# m1_11760_25858# pfet$348
Xpfet$360_4 vdd m1_33174_24224# m1_34278_25658# m1_32193_25858# pfet$360
Xpfet$350_26 vdd vdd vdd m1_16911_22102# m1_16452_21590# m1_16452_21590# pfet$350
Xpfet$350_15 vdd m1_354_22513# m1_354_22513# m1_n46_22402# m1_488_21786# m1_488_21786#
+ pfet$350
Xpfet$353_3 vdd vdd m1_n6657_17518# m1_n7247_17714# pfet$353
Xpfet$349_90 vdd m1_19747_15778# m1_18926_16202# m1_18665_17343# pfet$349
Xnfet$373_19 m1_n7513_20152# vss m1_1578_16080# vss nfet$373
Xpfet$351_0 vdd m1_2590_19404# m1_2590_19404# m1_3458_19550# m1_n3534_17714# m1_n3534_17714#
+ pfet$351
Xnfet$393_5 m1_26676_16080# m1_26676_16080# vss vss m1_28239_17358# vss nfet$393
Xnfet$379_3 m1_n1134_25662# m1_n290_24224# m1_814_25658# vss nfet$379
Xnfet$384_1 m1_28490_22513# m1_28490_22513# vss vss m1_34329_21430# vss nfet$384
Xnfet$377_0 m1_n3534_17714# vss m1_n6433_17343# vss nfet$377
Xpfet$376_2 vdd m1_n8283_20611# m1_n8283_20611# m1_n8047_22344# m1_n8145_21908# m1_n8145_21908#
+ pfet$376
Xpfet$369_1 vdd m1_n6856_24542# m1_n6856_24542# m1_n6624_23622# m1_n8283_19850# m1_n8283_19850#
+ pfet$369
Xnfet$370_7 m1_3049_25662# m1_3273_23922# m1_3537_24542# vss nfet$370
Xpfet$348_6 vdd vdd m1_3536_25662# m1_3394_25858# pfet$348
Xpfet$348_59 vdd vdd m1_16322_21786# pd6 pfet$348
Xpfet$348_48 vdd m1_16085_25662# m1_15822_23922# m1_15598_25662# pfet$348
Xpfet$348_37 vdd vdd m1_9973_24542# m1_7577_25858# pfet$348
Xpfet$348_26 vdd m1_4997_25658# m1_5790_24542# m1_3049_25662# pfet$348
Xpfet$348_15 vdd m1_11902_25662# m1_11639_23922# m1_11415_25662# pfet$348
Xpfet$360_5 vdd m1_32817_25662# m1_32554_23922# m1_32330_25662# pfet$360
Xpfet$350_27 vdd m1_14422_22513# m1_14422_22513# m1_14022_22402# m1_14556_21786# m1_14556_21786#
+ pfet$350
Xpfet$350_16 vdd m1_24973_22513# m1_24973_22513# m1_23945_22102# m1_25739_21786# m1_25739_21786#
+ pfet$350
Xpfet$353_4 vdd vdd m1_n6433_17343# m1_n3534_17714# pfet$353
Xpfet$349_91 vdd m1_24287_16080# m1_23820_18030# m1_22848_17343# pfet$349
Xpfet$349_80 vdd vdd m1_15564_15778# m1_15921_16080# pfet$349
Xpfet$351_1 vdd vdd vdd m1_2822_19850# m1_4620_20152# m1_4620_20152# pfet$351
Xnfet$379_4 m1_32193_25858# m1_34278_25658# m1_35071_24542# vss nfet$379
Xnfet$393_6 m1_27292_16202# m1_27292_16202# vss vss m1_26774_16398# vss nfet$393
Xnfet$384_2 m1_9645_21447# m1_9645_21447# vss vss m1_30492_21430# vss nfet$384
Xnfet$377_1 m1_n7513_20152# vss m1_n6788_16080# vss nfet$377
Xpfet$376_3 vdd vdd vdd m1_n8047_22344# m1_n8283_19850# m1_n8283_19850# pfet$376
Xpfet$348_7 vdd vdd m1_7232_25662# m1_7095_25858# pfet$348
Xnfet$370_8 m1_3394_25858# vss m1_3536_25662# vss nfet$370
Xpfet$348_49 vdd m1_20126_25858# vdd m1_21729_25658# pfet$348
Xpfet$348_38 vdd vdd m1_16085_25662# m1_15943_25858# pfet$348
Xpfet$348_27 vdd vdd m1_11278_25858# m1_7522_21786# pfet$348
Xpfet$348_16 vdd vdd m1_5771_21786# pd3 pfet$348
Xpfet$374_0 vdd vdd m1_n10796_25662# m1_n10933_25858# pfet$374
Xpfet$360_6 vdd m1_34278_25658# m1_35071_24542# m1_32330_25662# pfet$360
Xpfet$353_5 vdd vdd m1_n6788_16080# m1_n7513_20152# pfet$353
Xnfet$402_0 m1_n4485_21904# m1_n5764_21786# vss vss nfet$402
Xpfet$350_28 vdd m1_14422_22513# m1_14422_22513# m1_13394_22102# m1_15188_21786# m1_15188_21786#
+ pfet$350
Xpfet$350_17 vdd m1_21456_22513# m1_21456_22513# m1_21056_22402# m1_21590_21786# m1_21590_21786#
+ pfet$350
Xpfet$349_92 vdd m1_15454_18030# vdd m1_14127_16080# pfet$349
Xpfet$349_81 vdd vdd m1_13668_17714# m1_14127_16080# pfet$349
Xpfet$349_70 vdd vdd m1_18824_17836# m1_18665_17343# pfet$349
Xpfet$351_2 vdd m1_2590_19404# m1_2590_19404# m1_2822_19850# m1_2384_19550# m1_2384_19550#
+ pfet$351
Xnfet$379_5 m1_32330_25662# m1_33174_24224# m1_34278_25658# vss nfet$379
Xnfet$393_7 m1_26676_16080# m1_26676_16080# m1_26217_17714# m1_26217_17714# m1_26774_16398#
+ vss nfet$393
Xnfet$369_20 m1_21241_24346# m1_21241_24346# m1_20126_25858# m1_20126_25858# m1_22188_25502#
+ vss nfet$369
Xnfet$384_3 m1_7388_22513# m1_7388_22513# m1_30256_22102# m1_30256_22102# m1_30492_21430#
+ vss nfet$384
Xnfet$377_2 m1_n4994_16080# vss m1_n5351_15778# vss nfet$377
Xnfet$371_10 m1_19839_21786# m1_19839_21786# m1_21456_22513# m1_21456_22513# m1_21060_21586#
+ vss nfet$371
Xnfet$370_9 m1_3273_23922# vss m1_3893_24224# vss nfet$370
Xpfet$348_39 vdd vdd m1_15598_25662# m1_15461_25858# pfet$348
Xpfet$348_28 vdd m1_11639_23922# m1_11903_24542# m1_11278_25858# pfet$348
Xpfet$348_17 vdd vdd m1_7577_25858# m1_8692_24346# pfet$348
Xpfet$348_8 vdd vdd m1_8076_24224# m1_7456_23922# pfet$348
Xpfet$367_0 vdd m1_n4377_15778# m1_n4994_16080# m1_n6274_17836# pfet$367
Xpfet$374_1 vdd vdd m1_n10309_25662# m1_n10452_25858# pfet$374
Xnfet$382_0 m1_11039_21786# m1_11039_21786# vss vss m1_9877_21586# vss nfet$382
Xpfet$360_7 vdd m1_32554_23922# m1_32818_24542# m1_32193_25858# pfet$360
Xpfet$353_6 vdd vdd m1_n7383_17599# m1_n7247_17714# pfet$353
Xnfet$402_1 m1_n5227_21418# vss m1_n5764_21786# vss nfet$402
Xpfet$350_29 vdd vdd vdd m1_14022_22402# m1_12805_21786# m1_12805_21786# pfet$350
Xpfet$350_18 vdd vdd vdd m1_24573_22402# m1_23356_21786# m1_23356_21786# pfet$350
Xpfet$349_93 vdd m1_23820_18030# vdd m1_22493_16080# pfet$349
Xpfet$349_82 vdd m1_13668_17714# vdd m1_14743_16202# pfet$349
Xpfet$349_71 vdd vdd m1_19747_15778# m1_20104_16080# pfet$349
Xpfet$349_60 vdd vdd m1_n194_15778# m1_n3064_17714# pfet$349
Xpfet$351_3 vdd vdd vdd m1_3458_19550# m1_n3218_15478# m1_n3218_15478# pfet$351
Xnfet$374_10 m1_21590_21786# vss m1_22222_21786# vss nfet$374
Xnfet$379_6 m1_32193_25858# m1_32817_25662# m1_32554_23922# vss nfet$379
Xnfet$369_21 m1_28991_24224# m1_28991_24224# m1_28635_24542# m1_28635_24542# m1_29089_24542#
+ vss nfet$369
Xnfet$369_10 m1_17546_25658# m1_17546_25658# vss vss m1_18005_25502# vss nfet$369
Xnfet$377_3 m1_n6433_17343# vss m1_n6274_17836# vss nfet$377
Xnfet$371_11 m1_19969_21590# m1_19969_21590# m1_21456_22513# m1_21456_22513# m1_20428_21586#
+ vss nfet$371
Xnfet$382_10 m1_21590_21786# m1_21590_21786# vss vss m1_20428_21586# vss nfet$382
Xpfet$348_9 vdd m1_7719_25662# m1_7456_23922# m1_7232_25662# pfet$348
Xnfet$375_0 m1_n3534_17714# vss m1_2384_19550# vss nfet$375
Xnfet$382_1 m1_11671_21786# m1_11671_21786# vss vss m1_10509_21586# vss nfet$382
Xpfet$348_29 vdd vdd m1_11903_24542# m1_12259_24224# pfet$348
Xpfet$348_18 vdd vdd m1_11415_25662# m1_11278_25858# pfet$348
Xpfet$367_1 vdd m1_n5351_15778# m1_n6172_16202# m1_n6433_17343# pfet$367
Xpfet$374_2 vdd vdd m1_n9952_24224# m1_n10572_23922# pfet$374
Xpfet$353_7 vdd vdd m1_27190_17836# m1_27031_17343# pfet$353
Xnfet$402_2 m1_n6839_21786# vss m1_n6973_21481# vss nfet$402
Xpfet$350_19 vdd m1_24973_22513# m1_24973_22513# m1_24573_22402# m1_25107_21786# m1_25107_21786#
+ pfet$350
Xnfet$377_10 m1_26217_17714# vss m1_29087_15778# vss nfet$377
Xpfet$349_94 vdd vdd m1_22624_17518# m1_22034_17714# pfet$349
Xpfet$349_83 vdd m1_16538_15778# m1_15921_16080# m1_14641_17836# pfet$349
Xpfet$349_72 vdd m1_20721_15778# m1_20104_16080# m1_18824_17836# pfet$349
Xpfet$349_61 vdd m1_n811_16080# m1_n1278_18030# m1_n2250_17343# pfet$349
Xpfet$349_50 vdd m1_n1168_15778# m1_n1989_16202# m1_n2250_17343# pfet$349
Xpfet$351_4 vdd m1_6107_19404# m1_6107_19404# m1_6339_19850# m1_5901_19550# m1_5901_19550#
+ pfet$351
Xnfet$374_11 m1_18073_21786# vss m1_18705_21786# vss nfet$374
Xnfet$390_10 m1_9331_15478# m1_9331_15478# m1_n3822_21786# m1_n3822_21786# m1_13373_20470#
+ vss nfet$390
Xnfet$379_7 m1_32330_25662# m1_32554_23922# m1_32818_24542# vss nfet$379
Xnfet$369_22 m1_29607_24346# m1_29607_24346# vss vss m1_29089_24542# vss nfet$369
Xnfet$369_11 m1_16442_24224# m1_16442_24224# m1_16086_24542# m1_16086_24542# m1_16540_24542#
+ vss nfet$369
Xnfet$377_4 m1_n7247_17714# vss m1_n4377_15778# vss nfet$377
Xnfet$371_12 m1_16322_21786# m1_16322_21786# m1_17939_22513# m1_17939_22513# m1_17543_21586#
+ vss nfet$371
Xnfet$375_1 m1_n3218_15478# vss m1_4620_20152# vss nfet$375
Xnfet$382_2 m1_8154_21786# m1_8154_21786# vss vss m1_6992_21586# vss nfet$382
Xnfet$382_11 m1_22222_21786# m1_22222_21786# vss vss m1_21060_21586# vss nfet$382
Xpfet$348_19 vdd vdd m1_7095_25858# m1_4005_21786# pfet$348
Xpfet$367_2 vdd m1_n4994_16080# m1_n5461_18030# m1_n6433_17343# pfet$367
Xpfet$374_3 vdd vdd m1_n4978_24224# vss pfet$374
Xnfet$377_11 m1_27031_17343# vss m1_27190_17836# vss nfet$377
Xpfet$353_8 vdd vdd m1_28113_15778# m1_28470_16080# pfet$353
Xpfet$372_0 vdd vdd m1_n8625_26174# m1_n9336_24346# pfet$372
Xpfet$349_95 vdd vdd m1_21564_17714# m1_22034_17714# pfet$349
Xpfet$349_84 vdd vdd m1_17381_17714# m1_17851_17714# pfet$349
Xpfet$349_73 vdd vdd m1_16538_15778# m1_13668_17714# pfet$349
Xpfet$349_62 vdd vdd m1_23007_17836# m1_22848_17343# pfet$349
Xpfet$349_40 vdd m1_10560_16202# m1_10075_17518# m1_10458_17836# pfet$349
Xpfet$349_51 vdd vdd m1_n1168_15778# m1_n811_16080# pfet$349
Xpfet$351_5 vdd vdd vdd m1_n695_19850# m1_1103_20152# m1_1103_20152# pfet$351
Xnfet$400_0 m1_n7186_25858# vss m1_n7320_25516# vss nfet$400
Xpfet$351_30 vdd vdd vdd m1_24560_19550# m1_21880_15478# m1_21880_15478# pfet$351
Xnfet$374_12 m1_14556_21786# vss m1_15188_21786# vss nfet$374
Xnfet$390_11 m1_15171_20152# m1_15171_20152# m1_n3822_21786# m1_n3822_21786# m1_14005_20470#
+ vss nfet$390
Xnfet$369_23 m1_25424_24346# m1_25424_24346# m1_24309_25858# m1_24309_25858# m1_26371_25502#
+ vss nfet$369
Xnfet$369_12 m1_17058_24346# m1_17058_24346# m1_15943_25858# m1_15943_25858# m1_18005_25502#
+ vss nfet$369
Xnfet$398_0 m1_n9952_24224# m1_n9952_24224# m1_n10308_24542# m1_n10308_24542# m1_n9854_24542#
+ vss nfet$398
Xnfet$371_13 m1_16452_21590# m1_16452_21590# m1_17939_22513# m1_17939_22513# m1_16911_21586#
+ vss nfet$371
Xnfet$377_5 m1_n7247_17714# vss m1_n6657_17518# vss nfet$377
Xnfet$375_2 m1_n7401_15478# vss m1_1103_20152# vss nfet$375
Xnfet$382_3 m1_7522_21786# m1_7522_21786# vss vss m1_6360_21586# vss nfet$382
Xnfet$382_12 m1_18073_21786# m1_18073_21786# vss vss m1_16911_21586# vss nfet$382
Xpfet$367_3 vdd m1_n6172_16202# m1_n6657_17518# m1_n6274_17836# pfet$367
Xpfet$374_4 vdd vdd m1_n5571_25662# m1_n10452_25858# pfet$374
Xnfet$377_12 m1_28470_16080# vss m1_28113_15778# vss nfet$377
Xpfet$353_9 vdd vdd m1_29087_15778# m1_26217_17714# pfet$353
Xnfet$380_0 pd1 vss m1_n1263_21786# vss nfet$380
Xpfet$365_0 vdd m1_32818_20470# m1_32818_20470# m1_33050_19550# m1_30256_19792# m1_30256_19792#
+ pfet$365
Xpfet$372_1 vdd m1_n8625_26174# vdd m1_n8848_25658# pfet$372
Xpfet$349_96 vdd vdd m1_18665_17343# m1_21564_17714# pfet$349
Xpfet$349_85 vdd m1_18926_16202# m1_18441_17518# m1_18824_17836# pfet$349
Xpfet$349_74 vdd vdd m1_14641_17836# m1_14482_17343# pfet$349
Xpfet$349_63 vdd m1_23930_15778# m1_23109_16202# m1_22848_17343# pfet$349
Xpfet$349_30 vdd vdd m1_1933_17343# m1_4832_17714# pfet$349
Xpfet$349_41 vdd vdd m1_10075_17518# m1_9485_17714# pfet$349
Xpfet$349_52 vdd m1_n3064_17714# vdd m1_n1989_16202# pfet$349
Xnfet$400_1 m1_n6856_24542# vss m1_n6111_25858# vss nfet$400
Xpfet$351_6 vdd vdd vdd m1_6339_19850# m1_8137_20152# m1_8137_20152# pfet$351
Xpfet$351_31 vdd m1_n2543_20130# m1_n2543_20130# m1_20407_19850# m1_19969_19550# m1_19969_19550#
+ pfet$351
Xpfet$351_20 vdd m1_n3822_21786# m1_n3822_21786# m1_14009_19550# m1_9015_17714# m1_9015_17714#
+ pfet$351
Xnfet$374_13 m1_16322_21786# vss m1_16452_21590# vss nfet$374
Xnfet$390_12 m1_18688_20152# m1_18688_20152# m1_n1927_20274# m1_n1927_20274# m1_17522_20470#
+ vss nfet$390
Xnfet$369_24 m1_30095_25658# m1_30095_25658# vss vss m1_30554_25502# vss nfet$369
Xnfet$369_13 m1_13363_25658# m1_13363_25658# vss vss m1_13822_25502# vss nfet$369
Xnfet$398_1 m1_n9336_24346# m1_n9336_24346# m1_n8625_26174# m1_n8625_26174# m1_n8389_25502#
+ vss nfet$398
Xnfet$371_14 m1_12805_21786# m1_12805_21786# m1_14422_22513# m1_14422_22513# m1_14026_21586#
+ vss nfet$371
Xnfet$377_6 m1_n7247_17714# vss m1_n7383_17599# vss nfet$377
Xnfet$382_4 m1_1120_21786# m1_1120_21786# vss vss m1_n42_21586# vss nfet$382
Xnfet$382_13 m1_18705_21786# m1_18705_21786# vss vss m1_17543_21586# vss nfet$382
Xpfet$367_4 vdd m1_28113_15778# m1_27292_16202# m1_27031_17343# pfet$367
Xnfet$375_3 m1_649_17714# vss m1_5901_19550# vss nfet$375
Xpfet$374_5 vdd vdd m1_n4847_25662# m1_n10452_25858# pfet$374
Xnfet$377_13 m1_26217_17714# vss m1_25747_17714# vss nfet$377
Xnfet$380_1 pd2 vss m1_2254_21786# vss nfet$380
Xnfet$373_0 m1_9485_17714# vss m1_9015_17714# vss nfet$373
Xpfet$358_0 vdd vdd vdd m1_33050_22344# m1_31535_22102# m1_31535_22102# pfet$358
Xpfet$365_1 vdd vdd vdd m1_33050_19550# m1_31535_19792# m1_31535_19792# pfet$365
Xpfet$372_2 vdd m1_n3651_26174# vdd m1_n4978_24224# pfet$372
Xpfet$349_97 vdd vdd m1_22493_16080# m1_n7513_20152# pfet$349
Xpfet$349_86 vdd m1_19637_18030# vdd m1_18310_16080# pfet$349
Xpfet$349_75 vdd vdd m1_17697_15478# sd3 pfet$349
Xpfet$349_64 vdd vdd m1_23930_15778# m1_24287_16080# pfet$349
Xpfet$349_20 vdd vdd m1_1119_17714# m1_1578_16080# pfet$349
Xpfet$349_31 vdd m1_3372_16080# m1_2905_18030# m1_1933_17343# pfet$349
Xpfet$349_42 vdd m1_11271_18030# vdd m1_9944_16080# pfet$349
Xpfet$349_53 vdd vdd m1_n3218_15478# sd8 pfet$349
Xpfet$351_7 vdd vdd vdd m1_6975_19550# m1_965_15478# m1_965_15478# pfet$351
Xpfet$351_32 vdd m1_n2543_20130# m1_n2543_20130# m1_21043_19550# m1_17381_17714# m1_17381_17714#
+ pfet$351
Xpfet$351_21 vdd vdd vdd m1_13373_19850# m1_15171_20152# m1_15171_20152# pfet$351
Xpfet$351_10 vdd vdd vdd m1_9856_19850# m1_11654_20152# m1_11654_20152# pfet$351
Xnfet$374_14 m1_19839_21786# vss m1_19969_21590# vss nfet$374
Xnfet$390_13 m1_13514_15478# m1_13514_15478# m1_n1927_20274# m1_n1927_20274# m1_16890_20470#
+ vss nfet$390
Xnfet$369_25 m1_29607_24346# m1_29607_24346# m1_28492_25858# m1_28492_25858# m1_30554_25502#
+ vss nfet$369
Xnfet$369_14 m1_12875_24346# m1_12875_24346# m1_11760_25858# m1_11760_25858# m1_13822_25502#
+ vss nfet$369
Xnfet$398_2 m1_n8848_25658# m1_n8848_25658# vss vss m1_n8389_25502# vss nfet$398
Xnfet$377_7 m1_26217_17714# vss m1_26807_17518# vss nfet$377
Xnfet$371_15 m1_26873_21786# m1_26873_21786# m1_28490_22513# m1_28490_22513# m1_28094_21586#
+ vss nfet$371
Xpfet$349_110 vdd vdd m1_10458_17836# m1_10299_17343# pfet$349
Xnfet$382_14 m1_15188_21786# m1_15188_21786# vss vss m1_14026_21586# vss nfet$382
Xpfet$367_5 vdd m1_29087_15778# m1_28470_16080# m1_27190_17836# pfet$367
Xnfet$375_4 m1_4832_17714# vss m1_9418_19550# vss nfet$375
Xpfet$374_6 vdd vdd m1_n4623_25487# fin pfet$374
Xnfet$382_5 m1_4005_21786# m1_4005_21786# vss vss m1_2843_21586# vss nfet$382
Xnfet$380_2 pd9 vss m1_26873_21786# vss nfet$380
Xpfet$354_10 vdd vdd m1_29239_20152# m1_26063_15478# pfet$354
Xnfet$373_1 m1_9015_17714# vss m1_6116_17343# vss nfet$373
Xpfet$365_2 vdd m1_32818_21586# m1_32818_21586# m1_33050_22344# m1_30256_22102# m1_30256_22102#
+ pfet$365
Xpfet$372_3 vdd vdd m1_n3651_26174# m1_n3541_23922# pfet$372
Xpfet$349_98 vdd m1_20104_16080# m1_19637_18030# m1_18665_17343# pfet$349
Xpfet$349_87 vdd vdd m1_18310_16080# m1_n7513_20152# pfet$349
Xpfet$349_76 vdd m1_17851_17714# vdd m1_18926_16202# pfet$349
Xpfet$349_65 vdd m1_24904_15778# m1_24287_16080# m1_23007_17836# pfet$349
Xpfet$349_21 vdd vdd m1_965_15478# sd7 pfet$349
Xpfet$349_10 vdd m1_8172_15778# m1_7555_16080# m1_6275_17836# pfet$349
Xpfet$349_32 vdd vdd m1_2905_18030# m1_3015_15778# pfet$349
Xpfet$349_43 vdd vdd m1_11271_18030# m1_11381_15778# pfet$349
Xpfet$349_54 vdd vdd m1_n1278_18030# m1_n1168_15778# pfet$349
Xpfet$351_8 vdd m1_9624_19404# m1_9624_19404# m1_10492_19550# m1_4832_17714# m1_4832_17714#
+ pfet$351
Xpfet$351_33 vdd m1_n3206_20274# m1_n3206_20274# m1_24560_19550# m1_21564_17714# m1_21564_17714#
+ pfet$351
Xpfet$351_22 vdd vdd vdd m1_14009_19550# m1_9331_15478# m1_9331_15478# pfet$351
Xpfet$351_11 vdd vdd vdd m1_10492_19550# m1_5148_15478# m1_5148_15478# pfet$351
Xpfet$370_0 vdd m1_n10309_25662# m1_n10572_23922# m1_n10796_25662# pfet$370
Xnfet$374_15 m1_28624_21786# vss m1_29256_21786# vss nfet$374
Xnfet$390_14 m1_22205_20152# m1_22205_20152# m1_n2543_20130# m1_n2543_20130# m1_21039_20470#
+ vss nfet$390
Xnfet$398_3 m1_n9336_24346# m1_n9336_24346# vss vss m1_n9854_24542# vss nfet$398
Xnfet$369_26 m1_25912_25658# m1_25912_25658# vss vss m1_26371_25502# vss nfet$369
Xnfet$369_15 m1_25424_24346# m1_25424_24346# vss vss m1_24906_24542# vss nfet$369
Xnfet$377_8 m1_n7513_20152# vss m1_26676_16080# vss nfet$377
Xnfet$371_16 m1_27003_21590# m1_27003_21590# m1_28490_22513# m1_28490_22513# m1_27462_21586#
+ vss nfet$371
Xnfet$396_0 m1_n3822_20130# m1_n3822_20130# m1_n4485_20152# m1_n4485_20152# m1_n3724_20470#
+ vss nfet$396
Xpfet$349_100 vdd vdd m1_23820_18030# m1_23930_15778# pfet$349
Xnfet$382_15 m1_14556_21786# m1_14556_21786# vss vss m1_13394_21586# vss nfet$382
Xnfet$375_5 m1_965_15478# vss m1_8137_20152# vss nfet$375
Xnfet$382_6 m1_4637_21786# m1_4637_21786# vss vss m1_3475_21586# vss nfet$382
Xpfet$367_6 vdd m1_28470_16080# m1_28003_18030# m1_27031_17343# pfet$367
Xpfet$374_7 vdd vdd m1_n3541_23922# m1_n3184_24224# pfet$374
Xpfet$354_11 vdd vdd m1_18688_20152# m1_13514_15478# pfet$354
Xnfet$373_2 m1_6275_17836# m1_7555_16080# m1_7088_18030# vss nfet$373
Xpfet$372_4 vdd m1_n10452_25858# vdd m1_n4362_24346# pfet$372
Xpfet$349_99 vdd m1_23109_16202# m1_22624_17518# m1_23007_17836# pfet$349
Xpfet$349_88 vdd vdd m1_18441_17518# m1_17851_17714# pfet$349
Xpfet$349_77 vdd vdd m1_17851_17714# m1_18310_16080# pfet$349
Xpfet$349_66 vdd vdd m1_24904_15778# m1_22034_17714# pfet$349
Xpfet$349_22 vdd vdd m1_3015_15778# m1_3372_16080# pfet$349
Xpfet$349_11 vdd vdd m1_9485_17714# m1_9944_16080# pfet$349
Xpfet$349_33 vdd vdd m1_5892_17518# m1_5302_17714# pfet$349
Xpfet$349_44 vdd vdd m1_649_17714# m1_1119_17714# pfet$349
Xpfet$349_55 vdd vdd m1_n2474_17518# m1_n3064_17714# pfet$349
Xpfet$351_9 vdd m1_9624_19404# m1_9624_19404# m1_9856_19850# m1_9418_19550# m1_9418_19550#
+ pfet$351
Xpfet$363_0 vdd vdd vdd m1_36073_22344# define define pfet$363
Xpfet$351_34 vdd m1_n3206_20274# m1_n3206_20274# m1_23924_19850# m1_23486_19550# m1_23486_19550#
+ pfet$351
Xpfet$351_23 vdd vdd vdd m1_16890_19850# m1_18688_20152# m1_18688_20152# pfet$351
Xpfet$351_12 vdd m1_6107_19404# m1_6107_19404# m1_6975_19550# m1_649_17714# m1_649_17714#
+ pfet$351
Xpfet$370_1 vdd m1_n9952_24224# m1_n8848_25658# m1_n10933_25858# pfet$370
Xnfet$374_16 m1_26873_21786# vss m1_27003_21590# vss nfet$374
Xnfet$390_15 m1_17697_15478# m1_17697_15478# m1_n2543_20130# m1_n2543_20130# m1_20407_20470#
+ vss nfet$390
Xnfet$369_27 m1_12875_24346# m1_12875_24346# vss vss m1_12357_24542# vss nfet$369
Xnfet$369_16 m1_24808_24224# m1_24808_24224# m1_24452_24542# m1_24452_24542# m1_24906_24542#
+ vss nfet$369
Xnfet$398_4 m1_n4978_24224# m1_n4978_24224# m1_n10452_25858# m1_n10452_25858# m1_n4880_24542#
+ vss nfet$398
Xnfet$377_9 m1_n10452_25858# vss m1_27031_17343# vss nfet$377
Xnfet$371_17 m1_12935_21590# m1_12935_21590# m1_14422_22513# m1_14422_22513# m1_13394_21586#
+ vss nfet$371
Xnfet$389_0 m1_7198_15778# m1_7198_15778# m1_7088_18030# m1_7088_18030# m1_7324_17358#
+ vss nfet$389
Xnfet$396_1 m1_n1927_20274# m1_n1927_20274# vss vss m1_n2445_20470# vss nfet$396
Xpfet$349_101 vdd vdd m1_19637_18030# m1_19747_15778# pfet$349
Xnfet$382_7 m1_488_21786# m1_488_21786# vss vss m1_n674_21586# vss nfet$382
Xnfet$375_6 m1_9015_17714# vss m1_12935_19550# vss nfet$375
Xnfet$382_16 m1_28624_21786# m1_28624_21786# vss vss m1_27462_21586# vss nfet$382
Xpfet$367_7 vdd m1_27292_16202# m1_26807_17518# m1_27190_17836# pfet$367
Xpfet$374_8 vdd vdd m1_n2567_23922# m1_n7320_25516# pfet$374
Xpfet$354_12 vdd vdd m1_15171_20152# m1_9331_15478# pfet$354
Xnfet$373_3 m1_n7513_20152# vss m1_9944_16080# vss nfet$373
Xpfet$372_5 vdd vdd m1_n10308_24542# m1_n9952_24224# pfet$372
Xpfet$349_89 vdd vdd m1_22848_17343# m1_25747_17714# pfet$349
Xpfet$349_78 vdd vdd m1_13514_15478# sd4 pfet$349
Xpfet$349_67 vdd m1_22034_17714# vdd m1_23109_16202# pfet$349
Xpfet$349_12 vdd m1_3989_15778# m1_3372_16080# m1_2092_17836# pfet$349
Xpfet$349_23 vdd m1_5302_17714# vdd m1_6377_16202# pfet$349
Xpfet$349_34 vdd vdd m1_5761_16080# m1_n7513_20152# pfet$349
Xpfet$349_45 vdd vdd m1_9944_16080# m1_n7513_20152# pfet$349
Xpfet$349_56 vdd m1_n1278_18030# vdd m1_n2605_16080# pfet$349
Xnfet$371_0 m1_n1133_21590# m1_n1133_21590# m1_354_22513# m1_354_22513# m1_n674_21586#
+ vss nfet$371
Xpfet$363_1 vdd m1_35837_22102# m1_35837_22102# m1_36073_22344# fout fout pfet$363
Xpfet$370_2 vdd m1_n4362_24346# m1_n4847_25662# m1_n4464_25980# pfet$370
Xpfet$356_0 vdd vdd m1_n647_25662# m1_n789_25858# pfet$356
Xpfet$351_35 vdd m1_n3822_21786# m1_n3822_21786# m1_13373_19850# m1_12935_19550# m1_12935_19550#
+ pfet$351
Xpfet$351_24 vdd m1_n1927_20274# m1_n1927_20274# m1_16890_19850# m1_16452_19550# m1_16452_19550#
+ pfet$351
Xpfet$351_13 vdd m1_n927_19404# m1_n927_19404# m1_n695_19850# m1_n1133_19550# m1_n1133_19550#
+ pfet$351
Xnfet$374_17 m1_25107_21786# vss m1_25739_21786# vss nfet$374
Xnfet$390_16 m1_25722_20152# m1_25722_20152# m1_n3206_20274# m1_n3206_20274# m1_24556_20470#
+ vss nfet$390
Xnfet$369_17 m1_20625_24224# m1_20625_24224# m1_20269_24542# m1_20269_24542# m1_20723_24542#
+ vss nfet$369
Xnfet$398_5 m1_n4362_24346# m1_n4362_24346# vss vss m1_n4880_24542# vss nfet$398
Xnfet$389_1 m1_5761_16080# m1_5761_16080# vss vss m1_7324_17358# vss nfet$389
Xnfet$396_2 m1_n3206_20274# m1_n3206_20274# vss vss m1_n3724_20470# vss nfet$396
Xnfet$382_8 m1_25739_21786# m1_25739_21786# vss vss m1_24577_21586# vss nfet$382
Xpfet$349_102 vdd vdd m1_13198_17714# m1_13668_17714# pfet$349
Xnfet$375_7 m1_5148_15478# vss m1_11654_20152# vss nfet$375
Xnfet$382_17 m1_29256_21786# m1_29256_21786# vss vss m1_28094_21586# vss nfet$382
Xpfet$374_9 vdd vdd m1_n4464_25980# m1_n4623_25487# pfet$374
Xpfet$354_13 vdd vdd m1_16452_19550# m1_13198_17714# pfet$354
Xnfet$373_4 m1_10299_17343# m1_10560_16202# m1_10075_17518# vss nfet$373
Xpfet$349_13 vdd vdd m1_5148_15478# sd6 pfet$349
Xpfet$372_6 vdd m1_n10308_24542# vdd m1_n9336_24346# pfet$372
Xpfet$349_79 vdd m1_15564_15778# m1_14743_16202# m1_14482_17343# pfet$349
Xpfet$349_68 vdd vdd m1_22034_17714# m1_22493_16080# pfet$349
Xpfet$349_24 vdd m1_6377_16202# m1_5892_17518# m1_6275_17836# pfet$349
Xpfet$349_35 vdd vdd m1_9015_17714# m1_9485_17714# pfet$349
Xpfet$349_46 vdd vdd m1_n2250_17343# m1_649_17714# pfet$349
Xpfet$349_57 vdd m1_n1989_16202# m1_n2474_17518# m1_n2091_17836# pfet$349
Xpfet$349_0 vdd vdd m1_12355_15778# m1_9485_17714# pfet$349
Xnfet$371_1 m1_n1263_21786# m1_n1263_21786# m1_354_22513# m1_354_22513# m1_n42_21586#
+ vss nfet$371
Xpfet$356_1 vdd vdd m1_n1134_25662# m1_n1271_25858# pfet$356
Xpfet$370_3 vdd m1_n3184_24224# m1_n3651_26174# m1_n4623_25487# pfet$370
Xpfet$351_25 vdd vdd vdd m1_17526_19550# m1_13514_15478# m1_13514_15478# pfet$351
Xpfet$351_14 vdd m1_n927_19404# m1_n927_19404# m1_n59_19550# m1_n7383_17599# m1_n7383_17599#
+ pfet$351
Xnfet$390_17 m1_21880_15478# m1_21880_15478# m1_n3206_20274# m1_n3206_20274# m1_23924_20470#
+ vss nfet$390
Xnfet$369_18 m1_21241_24346# m1_21241_24346# vss vss m1_20723_24542# vss nfet$369
Xnfet$398_6 m1_n4978_24224# m1_n4978_24224# vss vss m1_n3415_25502# vss nfet$398
Xnfet$389_2 m1_9944_16080# m1_9944_16080# vss vss m1_11507_17358# vss nfet$389
Xnfet$396_3 m1_n6973_21481# m1_n6973_21481# m1_n6839_20152# m1_n6839_20152# m1_n6282_20470#
+ vss nfet$396
Xnfet$382_9 m1_25107_21786# m1_25107_21786# vss vss m1_23945_21586# vss nfet$382
Xpfet$349_103 vdd m1_14743_16202# m1_14258_17518# m1_14641_17836# pfet$349
Xnfet$375_8 m1_n7383_17599# vss m1_n1133_19550# vss nfet$375
Xnfet$394_0 m1_n10452_25858# m1_n10452_25858# m1_n7186_25858# m1_n7186_25858# m1_n6629_25502#
+ vss nfet$394
Xpfet$354_14 vdd vdd m1_23486_19550# m1_21564_17714# pfet$354
Xpfet$379_0 vdd vdd vdd m1_n5019_19550# m1_n4485_20152# m1_n4485_20152# pfet$379
Xnfet$373_5 m1_10458_17836# m1_11738_16080# m1_11271_18030# vss nfet$373
Xpfet$372_7 vdd vdd m1_n10452_25858# m1_n4978_24224# pfet$372
Xpfet$349_69 vdd vdd m1_20721_15778# m1_17851_17714# pfet$349
Xpfet$349_14 vdd vdd m1_2092_17836# m1_1933_17343# pfet$349
Xpfet$349_25 vdd vdd m1_1709_17518# m1_1119_17714# pfet$349
Xpfet$349_36 vdd vdd m1_6116_17343# m1_9015_17714# pfet$349
Xpfet$349_47 vdd m1_11738_16080# m1_11271_18030# m1_10299_17343# pfet$349
Xpfet$349_58 vdd vdd m1_n3534_17714# m1_n3064_17714# pfet$349
Xpfet$370_4 vdd m1_n2567_23922# m1_n3184_24224# m1_n4464_25980# pfet$370
Xnfet$371_2 m1_9288_21786# m1_9288_21786# m1_9645_21447# m1_9645_21447# m1_10509_21586#
+ vss nfet$371
Xpfet$351_26 vdd m1_n1927_20274# m1_n1927_20274# m1_17526_19550# m1_13198_17714# m1_13198_17714#
+ pfet$351
Xpfet$351_15 vdd vdd vdd m1_n59_19550# m1_n7401_15478# m1_n7401_15478# pfet$351
Xpfet$349_1 vdd vdd m1_11381_15778# m1_11738_16080# pfet$349
Xpfet$356_2 vdd vdd m1_n1271_25858# m1_n10452_25858# pfet$356
Xpfet$361_0 vdd vdd m1_n1263_21786# pd1 pfet$361
Xnfet$369_19 m1_21729_25658# m1_21729_25658# vss vss m1_22188_25502# vss nfet$369
Xnfet$398_7 m1_n3541_23922# m1_n3541_23922# m1_n3651_26174# m1_n3651_26174# m1_n3415_25502#
+ vss nfet$398
Xnfet$389_3 m1_11381_15778# m1_11381_15778# m1_11271_18030# m1_11271_18030# m1_11507_17358#
+ vss nfet$389
Xnfet$396_4 m1_2590_19404# m1_2590_19404# vss vss m1_n2445_21430# vss nfet$396
Xpfet$349_104 vdd vdd m1_14127_16080# m1_n7513_20152# pfet$349
Xnfet$375_9 m1_25747_17714# vss m1_27003_19550# vss nfet$375
Xnfet$394_1 m1_n6111_25858# m1_n6111_25858# vss vss m1_n6629_25502# vss nfet$394
Xnfet$387_0 m1_34093_22102# vss fout vss nfet$387
Xpfet$354_15 vdd vdd m1_22205_20152# m1_17697_15478# pfet$354
Xnfet$373_6 m1_6116_17343# vss m1_6275_17836# vss nfet$373
Xpfet$349_15 vdd vdd m1_5302_17714# m1_5761_16080# pfet$349
Xpfet$349_26 vdd vdd m1_4832_17714# m1_5302_17714# pfet$349
Xpfet$349_37 vdd m1_7555_16080# m1_7088_18030# m1_6116_17343# pfet$349
Xpfet$349_48 vdd vdd m1_n3064_17714# m1_n2605_16080# pfet$349
Xpfet$349_59 vdd vdd m1_n2605_16080# m1_n7513_20152# pfet$349
Xnfet$371_3 m1_9418_21590# m1_9418_21590# m1_9645_21447# m1_9645_21447# m1_9877_21586#
+ vss nfet$371
Xpfet$351_27 vdd vdd vdd m1_20407_19850# m1_22205_20152# m1_22205_20152# pfet$351
Xpfet$351_16 vdd vdd vdd m1_28077_19550# m1_26063_15478# m1_26063_15478# pfet$351
Xpfet$356_3 vdd vdd m1_1607_24542# m1_n789_25858# pfet$356
Xpfet$349_2 vdd m1_12355_15778# m1_11738_16080# m1_10458_17836# pfet$349
Xpfet$370_5 vdd m1_n10572_23922# m1_n10308_24542# m1_n10933_25858# pfet$370
Xpfet$361_1 vdd vdd m1_2254_21786# pd2 pfet$361
Xpfet$354_0 vdd vdd m1_2384_19550# m1_n3534_17714# pfet$354
Xnfet$389_4 m1_10560_16202# m1_10560_16202# vss vss m1_10042_16398# vss nfet$389
Xnfet$396_5 m1_6107_19404# m1_6107_19404# m1_n5227_21418# m1_n5227_21418# m1_n2445_21430#
+ vss nfet$396
Xpfet$349_105 vdd vdd m1_14258_17518# m1_13668_17714# pfet$349
Xpfet$354_16 vdd vdd m1_19969_19550# m1_17381_17714# pfet$354
Xnfet$373_7 m1_9485_17714# vss m1_10075_17518# vss nfet$373
Xpfet$349_16 vdd vdd m1_3989_15778# m1_1119_17714# pfet$349
Xpfet$349_27 vdd m1_2194_16202# m1_1709_17518# m1_2092_17836# pfet$349
Xpfet$349_38 vdd vdd m1_7088_18030# m1_7198_15778# pfet$349
Xpfet$349_49 vdd m1_n194_15778# m1_n811_16080# m1_n2091_17836# pfet$349
Xnfet$371_4 m1_5901_21590# m1_5901_21590# m1_7388_22513# m1_7388_22513# m1_6360_21586#
+ vss nfet$371
Xpfet$351_28 vdd vdd vdd m1_21043_19550# m1_17697_15478# m1_17697_15478# pfet$351
Xpfet$351_17 vdd m1_n3822_20130# m1_n3822_20130# m1_28077_19550# m1_25747_17714# m1_25747_17714#
+ pfet$351
Xpfet$356_4 vdd vdd m1_488_21786# m1_n789_25858# pfet$356
Xpfet$349_3 vdd m1_11381_15778# m1_10560_16202# m1_10299_17343# pfet$349
Xpfet$370_6 vdd m1_n8848_25658# m1_n8055_24542# m1_n10796_25662# pfet$370
Xpfet$361_2 vdd vdd m1_26873_21786# pd9 pfet$361
Xpfet$354_1 vdd vdd m1_4620_20152# m1_n3218_15478# pfet$354
Xnfet$389_5 m1_9944_16080# m1_9944_16080# m1_9485_17714# m1_9485_17714# m1_10042_16398#
+ vss nfet$389
Xnfet$396_6 m1_n5764_21786# m1_n5764_21786# vss vss m1_n6282_21430# vss nfet$396
Xpfet$349_106 vdd vdd m1_14482_17343# m1_17381_17714# pfet$349
Xpfet$354_17 vdd vdd m1_25722_20152# m1_21880_15478# pfet$354
Xnfet$372_10 m1_9015_17714# m1_9015_17714# vss vss m1_14005_20470# vss nfet$372
Xnfet$373_8 m1_7555_16080# vss m1_7198_15778# vss nfet$373
Xnfet$392_0 m1_n6274_17836# m1_n4994_16080# m1_n5461_18030# vss nfet$392
Xpfet$349_17 vdd vdd m1_n2091_17836# m1_n2250_17343# pfet$349
Xpfet$349_28 vdd m1_2905_18030# vdd m1_1578_16080# pfet$349
Xpfet$349_39 vdd m1_7088_18030# vdd m1_5761_16080# pfet$349
Xpfet$377_0 vdd m1_n6380_21786# m1_n6380_21786# m1_n5019_19550# m1_n5227_20152# m1_n5227_20152#
+ pfet$377
Xnfet$371_5 m1_2254_21786# m1_2254_21786# m1_3871_22513# m1_3871_22513# m1_3475_21586#
+ vss nfet$371
Xpfet$356_5 vdd vdd m1_326_24346# m1_n7513_20152# pfet$356
Xpfet$349_4 vdd m1_9485_17714# vdd m1_10560_16202# pfet$349
Xnfet$405_0 m1_n6839_20152# vss m1_n8145_21908# vss nfet$405
Xpfet$370_7 vdd m1_n3541_23922# m1_n4362_24346# m1_n4623_25487# pfet$370
Xpfet$351_29 vdd vdd vdd m1_23924_19850# m1_25722_20152# m1_25722_20152# pfet$351
Xpfet$351_18 vdd vdd vdd m1_27441_19850# m1_29239_20152# m1_29239_20152# pfet$351
Xpfet$354_2 vdd vdd m1_1103_20152# m1_n7401_15478# pfet$354
Xnfet$375_10 m1_26063_15478# vss m1_29239_20152# vss nfet$375
Xnfet$389_6 m1_1578_16080# m1_1578_16080# vss vss m1_3141_17358# vss nfet$389
Xnfet$396_7 m1_n3822_21786# m1_n3822_21786# m1_n4485_21904# m1_n4485_21904# m1_n3724_21430#
+ vss nfet$396
Xpfet$349_107 vdd m1_15921_16080# m1_15454_18030# m1_14482_17343# pfet$349
Xnfet$372_11 m1_13198_17714# m1_13198_17714# vss vss m1_17522_20470# vss nfet$372
Xnfet$373_9 sd5 vss m1_9331_15478# vss nfet$373
Xnfet$385_0 m1_31535_22102# m1_32818_21586# vss vss nfet$385
Xpfet$349_18 vdd m1_1119_17714# vdd m1_2194_16202# pfet$349
Xnfet$392_1 m1_n6433_17343# m1_n4377_15778# m1_n4994_16080# vss nfet$392
Xpfet$377_1 vdd vdd vdd m1_n5019_22344# m1_n4485_21904# m1_n4485_21904# pfet$377
Xpfet$349_29 vdd vdd m1_1578_16080# m1_n7513_20152# pfet$349
.ends

.subckt asc_drive_buffer$4 vss in vdd out
Xnfet$440_0 out out vss m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# m1_4274_n1060#
+ m1_4274_n1060# out m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# vss vss
+ nfet$440
Xpfet$416_0 vdd vdd m1_4002_n1060# m1_3466_n454# pfet$416
Xpfet$414_0 out out m1_4274_n1060# vdd m1_4274_n1060# out vdd vdd m1_4274_n1060# out
+ m1_4274_n1060# m1_4274_n1060# out m1_4274_n1060# vdd m1_4274_n1060# vdd m1_4274_n1060#
+ pfet$414
Xnfet$441_0 m1_3466_n454# vss m1_4002_n1060# vss nfet$441
Xpfet$417_0 vdd vdd m1_3466_n454# in pfet$417
Xpfet$415_0 m1_4274_n1060# vdd vdd m1_4274_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ vdd m1_4002_n1060# m1_4002_n1060# pfet$415
Xnfet$439_0 m1_4274_n1060# vss m1_4002_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ m1_4274_n1060# vss m1_4002_n1060# vss nfet$439
Xnfet$442_0 in vss m1_3466_n454# vss nfet$442
.ends

.subckt asc_hysteresis_buffer$8 vss in vdd out
Xpfet$389_0 vdd vdd m1_348_648# in pfet$389
Xpfet$387_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd
+ m1_884_42# m1_884_42# pfet$387
Xnfet$415_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$415
Xnfet$413_0 m1_348_648# vss m1_884_42# vss nfet$413
Xpfet$390_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$390
Xpfet$388_0 vdd vdd m1_884_42# m1_348_648# pfet$388
Xnfet$416_0 m1_1156_42# vss m1_884_42# vss nfet$416
Xnfet$414_0 in vss m1_348_648# vss nfet$414
Xpfet$391_0 vdd vdd m1_884_42# m1_1156_42# pfet$391
Xnfet$412_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$412
.ends

.subckt top_level_20250912_nosc$1 i_cp_100u div_def div_prc_s8 div_prc_s7 div_prc_s6
+ div_prc_s5 div_prc_s4 div_prc_s3 div_prc_s2 div_prc_s1 div_prc_s0 div_out div_in
+ div_swc_s0 div_swc_s1 div_swc_s2 div_swc_s3 div_swc_s4 div_swc_s5 div_swc_s6 div_swc_s7
+ div_swc_s8 ref ext_pfd_div ext_pfd_ref ext_pfd_up ext_pfd_down mx_pfd_s1 mx_pfd_s0
+ cp_s1 cp_s2 cp_s3 cp_s4 filter_in filter_out mx_vco_s0 mx_vco_s1 div_rpc_s0 div_rsc_s0
+ div_rsc_s1 div_rpc_s1 div_rsc_s2 div_rpc_s2 div_rsc_s3 div_rsc_s4 div_rsc_s5 div_rsc_s6
+ div_rsc_s7 div_rsc_s8 div_rpc_s3 div_rpc_s4 div_rpc_s5 div_rpc_s6 div_rpc_s7 div_rpc_s8
+ mx_ref_s1 mx_ref_s0 BIAS$2_0/200p1 BIAS$2_0/200n xp_3_1_MUX$4_0/B_1 xp_3_1_MUX$4_1/B_1
+ ext_vco_out up out down vdd lock ext_vco_in vss BIAS$2_0/200p2
Xxp_3_1_MUX$5_1 mx_ref_s0 mx_ref_s1 vdd vss xp_3_1_MUX$5_1/OUT_1 xp_3_1_MUX$5_1/C_1
+ xp_3_1_MUX$5_1/B_1 xp_3_1_MUX$5_1/A_1 xp_3_1_MUX$5
Xasc_dual_psd_def_20250809$5_0 vdd vss div_rpc_s0 div_rpc_s1 div_rpc_s2 div_rpc_s3
+ div_rpc_s4 div_rpc_s5 div_rpc_s6 div_rpc_s7 div_rpc_s8 xp_3_1_MUX$5_1/B_1 div_rsc_s0
+ div_rsc_s1 div_rsc_s2 div_rsc_s3 div_rsc_s4 div_rsc_s5 div_rsc_s6 div_rsc_s7 div_rsc_s8
+ xp_3_1_MUX$5_0/B_1 vss asc_dual_psd_def_20250809$5
Xasc_drive_buffer$5_0 vss xp_3_1_MUX$4_0/OUT_1 vdd asc_drive_buffer$4_0/in asc_drive_buffer$5
Xxp_programmable_basic_pump$2_0 asc_drive_buffer_up$2_0/out vdd cp_s1 cp_s2 cp_s3
+ cp_s4 asc_drive_buffer$4_6/out filter_in BIAS$2_0/100n vss xp_programmable_basic_pump$2
Xasc_PFD_DFF_20250831$2_0 vss xp_3_1_MUX$4_5/C_1 xp_3_1_MUX$4_2/C_1 vdd xp_3_1_MUX$4_4/C_1
+ xp_3_1_MUX$4_3/C_1 asc_PFD_DFF_20250831$2
Xasc_drive_buffer_up$2_0 vss asc_drive_buffer_up$2_0/out xp_3_1_MUX$4_2/OUT_1 vdd
+ asc_drive_buffer_up$2
Xasc_PFD_DFF_20250831$2_1 vss xp_3_1_MUX$4_2/B_1 xp_3_1_MUX$4_5/B_1 vdd xp_3_1_MUX$4_4/B_1
+ xp_3_1_MUX$4_3/B_1 asc_PFD_DFF_20250831$2
XBIAS$2_0 vdd vss BIAS$2_0/100n BIAS$2_0/200n i_cp_100u BIAS$2_0/200p1 BIAS$2_0/200p2
+ BIAS$2
Xasc_lock_detector_20250826$2_0 xp_3_1_MUX$4_3/OUT_1 vdd xp_3_1_MUX$4_4/OUT_1 vss
+ asc_drive_buffer$4_3/in asc_lock_detector_20250826$2
Xasc_hysteresis_buffer$7_0 vss xp_3_1_MUX$5_1/OUT_1 vdd xp_3_1_MUX$4_3/OUT_1 asc_hysteresis_buffer$7
XCSRVCO_20250823$2_0 xp_3_1_MUX$4_1/C_1 xp_3_1_MUX$4_0/C_1 vdd vss CSRVCO_20250823$2
Xxp_3_1_MUX$4_0 mx_vco_s0 mx_vco_s1 vdd vss xp_3_1_MUX$4_0/OUT_1 xp_3_1_MUX$4_0/C_1
+ xp_3_1_MUX$4_0/B_1 ext_vco_out xp_3_1_MUX$4
Xxp_3_1_MUX$4_1 mx_vco_s0 mx_vco_s1 vdd vss filter_out xp_3_1_MUX$4_1/C_1 xp_3_1_MUX$4_1/B_1
+ ext_vco_in xp_3_1_MUX$4
Xxp_3_1_MUX$4_2 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX$4_2/OUT_1 xp_3_1_MUX$4_2/C_1
+ xp_3_1_MUX$4_2/B_1 ext_pfd_up xp_3_1_MUX$4
Xxp_3_1_MUX$4_3 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX$4_3/OUT_1 xp_3_1_MUX$4_3/C_1
+ xp_3_1_MUX$4_3/B_1 ext_pfd_ref xp_3_1_MUX$4
Xasc_dual_psd_def_20250809$4_0 vdd vss div_prc_s0 div_prc_s1 div_prc_s2 div_prc_s3
+ div_prc_s4 div_prc_s5 div_prc_s6 div_prc_s7 div_prc_s8 xp_3_1_MUX$4_4/OUT_1 div_swc_s0
+ div_swc_s1 div_swc_s2 div_swc_s3 div_swc_s4 div_swc_s5 div_swc_s6 div_swc_s7 div_swc_s8
+ asc_drive_buffer$4_0/in div_def asc_dual_psd_def_20250809$4
Xxp_3_1_MUX$4_4 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX$4_4/OUT_1 xp_3_1_MUX$4_4/C_1
+ xp_3_1_MUX$4_4/B_1 ext_pfd_div xp_3_1_MUX$4
Xxp_3_1_MUX$4_5 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX$4_5/OUT_1 xp_3_1_MUX$4_5/C_1
+ xp_3_1_MUX$4_5/B_1 ext_pfd_down xp_3_1_MUX$4
Xasc_drive_buffer$4_1 vss xp_3_1_MUX$4_0/OUT_1 vdd out asc_drive_buffer$4
Xasc_drive_buffer$4_0 vss asc_drive_buffer$4_0/in vdd div_in asc_drive_buffer$4
Xasc_drive_buffer$4_2 vss xp_3_1_MUX$4_4/OUT_1 vdd div_out asc_drive_buffer$4
Xasc_drive_buffer$4_3 vss asc_drive_buffer$4_3/in vdd lock asc_drive_buffer$4
Xasc_drive_buffer$4_4 vss xp_3_1_MUX$4_2/OUT_1 vdd up asc_drive_buffer$4
Xasc_drive_buffer$4_5 vss xp_3_1_MUX$4_5/OUT_1 vdd down asc_drive_buffer$4
Xasc_drive_buffer$4_6 vss xp_3_1_MUX$4_5/OUT_1 vdd asc_drive_buffer$4_6/out asc_drive_buffer$4
Xasc_hysteresis_buffer$8_0 vss ref vdd xp_3_1_MUX$5_0/OUT_1 asc_hysteresis_buffer$8
Xxp_3_1_MUX$5_0 mx_ref_s0 mx_ref_s1 vdd vss xp_3_1_MUX$5_0/OUT_1 xp_3_1_MUX$5_1/C_1
+ xp_3_1_MUX$5_0/B_1 xp_3_1_MUX$5_0/A_1 xp_3_1_MUX$5
.ends

.subckt nfet$495 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$493 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$467 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$465 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$496 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$494 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$492 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$468 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$466 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$464 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt asc_hysteresis_buffer$10 vss vdd out in
Xnfet$495_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$495
Xnfet$493_0 m1_348_648# vss m1_884_42# vss nfet$493
Xpfet$467_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$467
Xpfet$465_0 vdd vdd m1_884_42# m1_348_648# pfet$465
Xnfet$496_0 m1_1156_42# vss m1_884_42# vss nfet$496
Xnfet$494_0 in vss m1_348_648# vss nfet$494
Xnfet$492_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$492
Xpfet$468_0 vdd vdd m1_884_42# m1_1156_42# pfet$468
Xpfet$466_0 vdd vdd m1_348_648# in pfet$466
Xpfet$464_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd
+ m1_884_42# m1_884_42# pfet$464
.ends

.subckt top_level_20250919_sc VDDd en clk ext_pfd_div ext_pfd_ref ext_pfd_down ext_pfd_up
+ i_cp_100u up filter_in filter_out out div_out data ref div_def ext_vco_out down
+ lock ext_vco_in div_in VSSd
Xscan_chain$1_0 VDDd en data clk scan_chain$1_0/out[1] scan_chain$1_0/out[2] scan_chain$1_0/out[3]
+ scan_chain$1_0/out[4] scan_chain$1_0/out[5] scan_chain$1_0/out[6] scan_chain$1_0/out[7]
+ scan_chain$1_0/out[8] scan_chain$1_0/out[9] scan_chain$1_0/out[10] scan_chain$1_0/out[20]
+ scan_chain$1_0/out[19] scan_chain$1_0/out[18] scan_chain$1_0/out[17] scan_chain$1_0/out[16]
+ scan_chain$1_0/out[15] scan_chain$1_0/out[14] scan_chain$1_0/out[13] scan_chain$1_0/out[12]
+ scan_chain$1_0/out[11] scan_chain$1_0/out[21] scan_chain$1_0/out[22] scan_chain$1_0/out[23]
+ scan_chain$1_0/out[24] scan_chain$1_0/out[25] scan_chain$1_0/out[26] VCOfinal$1_0/s0
+ VCOfinal$1_0/s1 VCOfinal$1_0/s2 VCOfinal$1_0/s3 scan_chain$1_0/out[40] scan_chain$1_0/out[39]
+ scan_chain$1_0/out[38] scan_chain$1_0/out[37] scan_chain$1_0/out[36] scan_chain$1_0/out[35]
+ scan_chain$1_0/out[34] scan_chain$1_0/out[33] scan_chain$1_0/out[32] scan_chain$1_0/out[31]
+ scan_chain$1_0/out[41] scan_chain$1_0/out[42] scan_chain$1_0/out[43] scan_chain$1_0/out[44]
+ scan_chain$1_0/out[45] scan_chain$1_0/out[46] scan_chain$1_0/out[47] scan_chain$1_0/out[48]
+ scan_chain$1_0/out[49] scan_chain$1_0/out[50] VSSd scan_chain$1
XVCOfinal$1_0 VCOfinal$1_0/s3 VCOfinal$1_0/s0 VCOfinal$1_0/s1 VCOfinal$1_0/s2 VCOfinal$1_0/iref200
+ VCOfinal$1_0/fout VCOfinal$1_0/foutb VCOfinal$1_0/irefp VCOfinal$1_0/irefn VCOfinal$1_0/vin
+ VSSd VDDd VSSd VCOfinal$1
Xtop_level_20250912_nosc$1_0 i_cp_100u asc_hysteresis_buffer$10_0/out scan_chain$1_0/out[42]
+ scan_chain$1_0/out[43] scan_chain$1_0/out[44] scan_chain$1_0/out[45] scan_chain$1_0/out[46]
+ scan_chain$1_0/out[47] scan_chain$1_0/out[48] scan_chain$1_0/out[49] scan_chain$1_0/out[50]
+ div_out div_in scan_chain$1_0/out[41] scan_chain$1_0/out[40] scan_chain$1_0/out[39]
+ scan_chain$1_0/out[38] scan_chain$1_0/out[37] scan_chain$1_0/out[36] scan_chain$1_0/out[35]
+ scan_chain$1_0/out[34] scan_chain$1_0/out[33] ref ext_pfd_div ext_pfd_ref ext_pfd_up
+ ext_pfd_down scan_chain$1_0/out[1] scan_chain$1_0/out[2] scan_chain$1_0/out[6] scan_chain$1_0/out[5]
+ scan_chain$1_0/out[4] scan_chain$1_0/out[3] filter_in filter_out scan_chain$1_0/out[32]
+ scan_chain$1_0/out[31] scan_chain$1_0/out[26] scan_chain$1_0/out[17] scan_chain$1_0/out[16]
+ scan_chain$1_0/out[25] scan_chain$1_0/out[15] scan_chain$1_0/out[24] scan_chain$1_0/out[14]
+ scan_chain$1_0/out[13] scan_chain$1_0/out[12] scan_chain$1_0/out[11] scan_chain$1_0/out[10]
+ scan_chain$1_0/out[9] scan_chain$1_0/out[23] scan_chain$1_0/out[22] scan_chain$1_0/out[21]
+ scan_chain$1_0/out[20] scan_chain$1_0/out[19] scan_chain$1_0/out[18] scan_chain$1_0/out[7]
+ scan_chain$1_0/out[8] VCOfinal$1_0/iref200 VCOfinal$1_0/irefn VCOfinal$1_0/fout
+ VCOfinal$1_0/vin ext_vco_out up out down VDDd lock ext_vco_in VSSd VCOfinal$1_0/irefp
+ top_level_20250912_nosc$1
Xasc_hysteresis_buffer$10_0 VSSd VDDd asc_hysteresis_buffer$10_0/out div_def asc_hysteresis_buffer$10
.ends

.subckt top_level_20250921 ref ext_pfd_div ext_pfd_ref ext_pfd_up ext_pfd_down lock
+ i_cp_100u up filter_in ext_vco_out ext_vco_in filter_out out div_in div_out div_def
+ clk data en VSSd VDDd down
XDECAP_LARGE_0 VDDd VSSd DECAP_LARGE
Xppolyf_u_resistor$9_0 VSSd top_level_20250919_sc_0/en VSSd ppolyf_u_resistor$9
Xio_secondary_3p3_0 data VDDd VSSd io_secondary_3p3_0/to_gate io_secondary_3p3
Xio_secondary_3p3_1 en VDDd VSSd top_level_20250919_sc_0/en io_secondary_3p3
Xio_secondary_3p3_2 div_def VDDd VSSd io_secondary_3p3_2/to_gate io_secondary_3p3
Xio_secondary_3p3_4 ref VDDd VSSd io_secondary_3p3_4/to_gate io_secondary_3p3
Xppolyf_u_resistor_0 VSSd ext_pfd_div top_level_20250919_sc_0/ext_pfd_div ppolyf_u_resistor
Xio_secondary_3p3_3 clk VDDd VSSd io_secondary_3p3_3/to_gate io_secondary_3p3
Xio_secondary_3p3_5 i_cp_100u VDDd VSSd io_secondary_3p3_5/to_gate io_secondary_3p3
Xppolyf_u_resistor_1 VSSd ext_pfd_up top_level_20250919_sc_0/ext_pfd_up ppolyf_u_resistor
Xppolyf_u_resistor_2 VSSd ext_pfd_ref top_level_20250919_sc_0/ext_pfd_ref ppolyf_u_resistor
Xppolyf_u_resistor_3 VSSd div_in top_level_20250919_sc_0/div_in ppolyf_u_resistor
Xtop_level_20250919_sc_0 VDDd top_level_20250919_sc_0/en io_secondary_3p3_3/to_gate
+ top_level_20250919_sc_0/ext_pfd_div top_level_20250919_sc_0/ext_pfd_ref top_level_20250919_sc_0/ext_pfd_down
+ top_level_20250919_sc_0/ext_pfd_up io_secondary_3p3_5/to_gate top_level_20250919_sc_0/up
+ top_level_20250919_sc_0/filter_in top_level_20250919_sc_0/filter_out top_level_20250919_sc_0/out
+ top_level_20250919_sc_0/div_out io_secondary_3p3_0/to_gate io_secondary_3p3_4/to_gate
+ io_secondary_3p3_2/to_gate top_level_20250919_sc_0/ext_vco_out top_level_20250919_sc_0/down
+ top_level_20250919_sc_0/lock top_level_20250919_sc_0/ext_vco_in top_level_20250919_sc_0/div_in
+ VSSd top_level_20250919_sc
Xppolyf_u_resistor_4 VSSd out top_level_20250919_sc_0/out ppolyf_u_resistor
Xppolyf_u_resistor_5 VSSd filter_out top_level_20250919_sc_0/filter_out ppolyf_u_resistor
Xppolyf_u_resistor_6 VSSd ext_vco_in top_level_20250919_sc_0/ext_vco_in ppolyf_u_resistor
Xppolyf_u_resistor_7 VSSd ext_vco_out top_level_20250919_sc_0/ext_vco_out ppolyf_u_resistor
Xppolyf_u_resistor_10 VSSd up top_level_20250919_sc_0/up ppolyf_u_resistor
Xppolyf_u_resistor_8 VSSd filter_in top_level_20250919_sc_0/filter_in ppolyf_u_resistor
Xppolyf_u_resistor_11 VSSd lock top_level_20250919_sc_0/lock ppolyf_u_resistor
Xppolyf_u_resistor_9 VSSd down top_level_20250919_sc_0/down ppolyf_u_resistor
Xppolyf_u_resistor_12 VSSd div_out top_level_20250919_sc_0/div_out ppolyf_u_resistor
Xppolyf_u_resistor_13 VSSd ext_pfd_down top_level_20250919_sc_0/ext_pfd_down ppolyf_u_resistor
.ends

