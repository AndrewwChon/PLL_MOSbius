* NGSPICE file created from top_level_20250919_sc.ext - technology: gf180mcuD

.subckt pfet$203 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$201 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$218 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$216 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt nfet$214 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$204 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$202 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$217 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$215 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$205 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt asc_drive_buffer_up vss out in vdd
Xpfet$203_0 vdd vdd m1_506_712# m1_n30_1318# pfet$203
Xpfet$201_0 out out m1_778_712# vdd m1_778_712# out vdd vdd m1_778_712# out m1_778_712#
+ m1_778_712# out m1_778_712# vdd m1_778_712# vdd m1_778_712# pfet$201
Xnfet$218_0 in vss m1_n566_1318# vss nfet$218
Xnfet$216_0 m1_n30_1318# vss m1_506_712# vss nfet$216
Xnfet$214_0 m1_778_712# vss m1_506_712# m1_506_712# m1_506_712# m1_778_712# m1_778_712#
+ vss m1_506_712# vss nfet$214
Xpfet$204_0 vdd vdd m1_n30_1318# m1_n566_1318# pfet$204
Xpfet$202_0 m1_778_712# vdd vdd m1_778_712# m1_506_712# m1_506_712# m1_778_712# vdd
+ m1_506_712# m1_506_712# pfet$202
Xnfet$217_0 m1_n566_1318# vss m1_n30_1318# vss nfet$217
Xnfet$215_0 out out vss m1_778_712# m1_778_712# out vss m1_778_712# m1_778_712# m1_778_712#
+ out m1_778_712# m1_778_712# out vss m1_778_712# vss vss nfet$215
Xpfet$205_0 vdd vdd m1_n566_1318# in pfet$205
.ends

.subckt nfet$169 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$159 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$166 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$154 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$170 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$172 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$158 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$142 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$164 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$149 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$151 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$155 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$163 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$162 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$148 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$141 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$162 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$145 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$156 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$160 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$153 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$179 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$161 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$146 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$140 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$184 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$169 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$151 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$177 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$152 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$144 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$155 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$182 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$167 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$175 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$168 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$143 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$172 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$150 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$180 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$165 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$153 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$173 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$158 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$166 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$170 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$159 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$163 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$156 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$171 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$164 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$149 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$157 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$161 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$154 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$147 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$185 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$152 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$178 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$160 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$183 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$168 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$150 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$176 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$181 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$174 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$167 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$171 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$157 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$165 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_dual_psd_def_20250809 vdd vss pd1 pd2 pd3 pd4 pd5 pd6 pd7 pd8 pd9 fout
+ sd1 sd2 sd3 sd4 sd5 sd6 sd7 sd8 sd9 fin define
Xnfet$169_9 m1_2194_16202# m1_2194_16202# vss vss m1_1676_16398# vss nfet$169
Xpfet$159_7 vdd m1_27292_16202# m1_26807_17518# m1_27190_17836# pfet$159
Xpfet$166_8 vdd vdd m1_n2567_23922# m1_n7320_25516# pfet$166
Xnfet$154_15 m1_28624_21786# vss m1_29256_21786# vss nfet$154
Xnfet$170_14 m1_22205_20152# m1_22205_20152# m1_n2543_20130# m1_n2543_20130# m1_21039_20470#
+ vss nfet$170
Xnfet$172_4 m1_27031_17343# m1_27292_16202# m1_26807_17518# vss nfet$172
Xnfet$158_2 m1_n1271_25858# vss m1_n1134_25662# vss nfet$158
Xpfet$142_32 vdd m1_28490_22513# m1_28490_22513# m1_28090_22402# m1_28624_21786# m1_28624_21786#
+ pfet$142
Xpfet$142_21 vdd vdd vdd m1_21056_22402# m1_19839_21786# m1_19839_21786# pfet$142
Xpfet$164_5 vdd vdd m1_n10308_24542# m1_n9952_24224# pfet$164
Xpfet$142_10 vdd m1_3871_22513# m1_3871_22513# m1_2843_22102# m1_4637_21786# m1_4637_21786#
+ pfet$142
Xnfet$149_26 m1_25912_25658# m1_25912_25658# vss vss m1_26371_25502# vss nfet$149
Xnfet$149_15 m1_25424_24346# m1_25424_24346# vss vss m1_24906_24542# vss nfet$149
Xnfet$151_9 m1_23356_21786# m1_23356_21786# m1_24973_22513# m1_24973_22513# m1_24577_21586#
+ vss nfet$151
Xnfet$170_1 m1_1103_20152# m1_1103_20152# m1_n927_19404# m1_n927_19404# m1_n63_20470#
+ vss nfet$170
Xpfet$155_1 vdd m1_35837_22102# m1_35837_22102# m1_36073_22344# fout fout pfet$155
Xnfet$163_0 m1_21456_22513# m1_21456_22513# m1_30256_19792# m1_30256_19792# m1_30492_20470#
+ vss nfet$163
Xpfet$162_2 vdd m1_n4362_24346# m1_n4847_25662# m1_n4464_25980# pfet$162
Xpfet$148_0 vdd vdd m1_n647_25662# m1_n789_25858# pfet$148
Xnfet$151_16 m1_27003_21590# m1_27003_21590# m1_28490_22513# m1_28490_22513# m1_27462_21586#
+ vss nfet$151
Xpfet$141_7 vdd vdd m1_6275_17836# m1_6116_17343# pfet$141
Xnfet$162_15 m1_14556_21786# m1_14556_21786# vss vss m1_13394_21586# vss nfet$162
Xpfet$145_10 vdd vdd m1_27031_17343# m1_n10452_25858# pfet$145
Xpfet$166_9 vdd vdd m1_n4464_25980# m1_n4623_25487# pfet$166
Xnfet$154_16 m1_26873_21786# vss m1_27003_21590# vss nfet$154
Xnfet$170_15 m1_17697_15478# m1_17697_15478# m1_n2543_20130# m1_n2543_20130# m1_20407_20470#
+ vss nfet$170
Xnfet$172_5 m1_27031_17343# m1_29087_15778# m1_28470_16080# vss nfet$172
Xnfet$158_3 m1_n7513_20152# vss m1_326_24346# vss nfet$158
Xpfet$142_33 vdd m1_28490_22513# m1_28490_22513# m1_27462_22102# m1_29256_21786# m1_29256_21786#
+ pfet$142
Xpfet$142_22 vdd m1_21456_22513# m1_21456_22513# m1_20428_22102# m1_22222_21786# m1_22222_21786#
+ pfet$142
Xpfet$164_6 vdd m1_n10308_24542# vdd m1_n9336_24346# pfet$164
Xpfet$142_11 vdd vdd vdd m1_2843_22102# m1_2384_21590# m1_2384_21590# pfet$142
Xnfet$149_27 m1_12875_24346# m1_12875_24346# vss vss m1_12357_24542# vss nfet$149
Xnfet$149_16 m1_24808_24224# m1_24808_24224# m1_24452_24542# m1_24452_24542# m1_24906_24542#
+ vss nfet$149
Xnfet$163_1 m1_14422_22513# m1_14422_22513# m1_31535_19792# m1_31535_19792# m1_31771_20470#
+ vss nfet$163
Xnfet$170_2 m1_n3218_15478# m1_n3218_15478# m1_2590_19404# m1_2590_19404# m1_2822_20470#
+ vss nfet$170
Xnfet$156_0 sd9 vss m1_n7401_15478# vss nfet$156
Xpfet$162_3 vdd m1_n3184_24224# m1_n3651_26174# m1_n4623_25487# pfet$162
Xnfet$151_17 m1_12935_21590# m1_12935_21590# m1_14422_22513# m1_14422_22513# m1_13394_21586#
+ vss nfet$151
Xpfet$148_1 vdd vdd m1_n1134_25662# m1_n1271_25858# pfet$148
Xpfet$141_8 vdd vdd m1_9331_15478# sd5 pfet$141
Xpfet$148_10 vdd vdd m1_35071_24542# m1_32675_25947# pfet$148
Xpfet$160_0 vdd vdd m1_n7513_20152# m1_35837_22102# pfet$160
Xnfet$162_16 m1_28624_21786# m1_28624_21786# vss vss m1_27462_21586# vss nfet$162
Xpfet$145_11 vdd vdd m1_26807_17518# m1_26217_17714# pfet$145
Xnfet$154_17 m1_25107_21786# vss m1_25739_21786# vss nfet$154
Xnfet$170_16 m1_25722_20152# m1_25722_20152# m1_n3206_20274# m1_n3206_20274# m1_24556_20470#
+ vss nfet$170
Xnfet$172_6 m1_27190_17836# m1_28113_15778# m1_27292_16202# vss nfet$172
Xnfet$158_4 m1_n789_25858# vss m1_1607_24542# vss nfet$158
Xpfet$142_34 vdd vdd vdd m1_28090_22402# m1_26873_21786# m1_26873_21786# pfet$142
Xpfet$142_23 vdd vdd vdd m1_23945_22102# m1_23486_21590# m1_23486_21590# pfet$142
Xpfet$164_7 vdd vdd m1_n10452_25858# m1_n4978_24224# pfet$164
Xpfet$142_12 vdd vdd vdd m1_3471_22402# m1_2254_21786# m1_2254_21786# pfet$142
Xnfet$149_17 m1_20625_24224# m1_20625_24224# m1_20269_24542# m1_20269_24542# m1_20723_24542#
+ vss nfet$149
Xnfet$156_1 sd2 vss m1_21880_15478# vss nfet$156
Xnfet$163_2 m1_17939_22513# m1_17939_22513# vss vss m1_31771_20470# vss nfet$163
Xnfet$170_3 m1_8137_20152# m1_8137_20152# m1_6107_19404# m1_6107_19404# m1_6971_20470#
+ vss nfet$170
Xnfet$149_0 m1_4509_24346# m1_4509_24346# vss vss m1_3991_24542# vss nfet$149
Xpfet$162_4 vdd m1_n2567_23922# m1_n3184_24224# m1_n4464_25980# pfet$162
Xpfet$148_2 vdd vdd m1_n1271_25858# m1_n10452_25858# pfet$148
Xpfet$141_9 vdd vdd m1_8172_15778# m1_5302_17714# pfet$141
Xpfet$148_11 vdd vdd m1_32817_25662# m1_32675_25947# pfet$148
Xpfet$153_0 vdd vdd m1_n1263_21786# pd1 pfet$153
Xnfet$162_17 m1_29256_21786# m1_29256_21786# vss vss m1_28094_21586# vss nfet$162
Xpfet$145_12 vdd vdd m1_26676_16080# m1_n7513_20152# pfet$145
Xnfet$179_0 m1_n10933_25858# m1_n8848_25658# m1_n8055_24542# vss nfet$179
Xnfet$170_17 m1_21880_15478# m1_21880_15478# m1_n3206_20274# m1_n3206_20274# m1_23924_20470#
+ vss nfet$170
Xnfet$172_7 m1_27190_17836# m1_28470_16080# m1_28003_18030# vss nfet$172
Xnfet$158_5 m1_n789_25858# vss m1_488_21786# vss nfet$158
Xpfet$142_35 vdd vdd vdd m1_13394_22102# m1_12935_21590# m1_12935_21590# pfet$142
Xnfet$149_18 m1_21241_24346# m1_21241_24346# vss vss m1_20723_24542# vss nfet$149
Xpfet$142_24 vdd m1_17939_22513# m1_17939_22513# m1_16911_22102# m1_18705_21786# m1_18705_21786#
+ pfet$142
Xpfet$142_13 vdd vdd vdd m1_6988_22402# m1_5771_21786# m1_5771_21786# pfet$142
Xnfet$156_2 sd1 vss m1_26063_15478# vss nfet$156
Xnfet$163_3 m1_24973_22513# m1_24973_22513# vss vss m1_30492_20470# vss nfet$163
Xnfet$170_4 m1_965_15478# m1_965_15478# m1_6107_19404# m1_6107_19404# m1_6339_20470#
+ vss nfet$170
Xnfet$149_1 m1_3893_24224# m1_3893_24224# m1_3537_24542# m1_3537_24542# m1_3991_24542#
+ vss nfet$149
Xpfet$148_3 vdd vdd m1_1607_24542# m1_n789_25858# pfet$148
Xpfet$162_5 vdd m1_n10572_23922# m1_n10308_24542# m1_n10933_25858# pfet$162
Xpfet$148_12 vdd vdd m1_32193_25858# m1_25107_21786# pfet$148
Xnfet$161_0 m1_n290_24224# m1_n290_24224# m1_n646_24542# m1_n646_24542# m1_n192_24542#
+ vss nfet$161
Xpfet$153_1 vdd vdd m1_2254_21786# pd2 pfet$153
Xpfet$146_0 vdd vdd m1_2384_19550# m1_n3534_17714# pfet$146
Xpfet$140_90 vdd vdd m1_24309_25858# m1_25424_24346# pfet$140
Xpfet$145_13 vdd vdd m1_25747_17714# m1_26217_17714# pfet$145
Xnfet$179_1 m1_n10796_25662# m1_n10572_23922# m1_n10308_24542# vss nfet$179
Xnfet$158_6 m1_n910_23922# vss m1_n290_24224# vss nfet$158
Xnfet$149_19 m1_21729_25658# m1_21729_25658# vss vss m1_22188_25502# vss nfet$149
Xpfet$142_25 vdd m1_17939_22513# m1_17939_22513# m1_17539_22402# m1_18073_21786# m1_18073_21786#
+ pfet$142
Xpfet$142_14 vdd vdd vdd m1_n46_22402# m1_n1263_21786# m1_n1263_21786# pfet$142
Xnfet$163_4 m1_32818_20470# m1_32818_20470# vss vss m1_34329_20470# vss nfet$163
Xnfet$149_2 m1_4997_25658# m1_4997_25658# vss vss m1_5456_25502# vss nfet$149
Xnfet$170_5 m1_5148_15478# m1_5148_15478# m1_9624_19404# m1_9624_19404# m1_9856_20470#
+ vss nfet$170
Xpfet$148_4 vdd vdd m1_488_21786# m1_n789_25858# pfet$148
Xpfet$162_6 vdd m1_n8848_25658# m1_n8055_24542# m1_n10796_25662# pfet$162
Xnfet$161_1 m1_814_25658# m1_814_25658# vss vss m1_1273_25502# vss nfet$161
Xnfet$154_0 m1_n1263_21786# vss m1_n1133_21590# vss nfet$154
Xpfet$148_13 vdd vdd m1_33790_24346# m1_n7513_20152# pfet$148
Xpfet$153_2 vdd vdd m1_26873_21786# pd9 pfet$153
Xpfet$146_1 vdd vdd m1_4620_20152# m1_n3218_15478# pfet$146
Xpfet$140_91 vdd vdd m1_23356_21786# pd8 pfet$140
Xpfet$140_80 vdd vdd m1_17058_24346# m1_n7513_20152# pfet$140
Xnfet$179_2 m1_n10933_25858# m1_n10309_25662# m1_n10572_23922# vss nfet$179
Xnfet$158_7 m1_25107_21786# vss m1_32193_25858# vss nfet$158
Xpfet$142_26 vdd vdd vdd m1_16911_22102# m1_16452_21590# m1_16452_21590# pfet$142
Xpfet$142_15 vdd m1_354_22513# m1_354_22513# m1_n46_22402# m1_488_21786# m1_488_21786#
+ pfet$142
Xnfet$184_0 m1_n4485_20152# m1_n6380_21786# vss vss nfet$184
Xpfet$169_0 vdd m1_n6380_21786# m1_n6380_21786# m1_n5019_19550# m1_n5227_20152# m1_n5227_20152#
+ pfet$169
Xnfet$170_6 m1_11654_20152# m1_11654_20152# m1_9624_19404# m1_9624_19404# m1_10488_20470#
+ vss nfet$170
Xnfet$163_5 m1_32818_21586# m1_32818_21586# m1_34093_19792# m1_34093_19792# m1_34329_20470#
+ vss nfet$163
Xpfet$148_5 vdd vdd m1_326_24346# m1_n7513_20152# pfet$148
Xnfet$149_3 m1_4509_24346# m1_4509_24346# m1_3394_25858# m1_3394_25858# m1_5456_25502#
+ vss nfet$149
Xpfet$162_7 vdd m1_n3541_23922# m1_n4362_24346# m1_n4623_25487# pfet$162
Xnfet$161_2 m1_326_24346# m1_326_24346# m1_n789_25858# m1_n789_25858# m1_1273_25502#
+ vss nfet$161
Xnfet$154_1 m1_11039_21786# vss m1_11671_21786# vss nfet$154
Xpfet$146_2 vdd vdd m1_1103_20152# m1_n7401_15478# pfet$146
Xpfet$140_92 vdd vdd m1_28492_25858# m1_29607_24346# pfet$140
Xpfet$140_81 vdd vdd m1_18339_24542# m1_15943_25858# pfet$140
Xpfet$140_70 vdd vdd m1_14156_24542# m1_11760_25858# pfet$140
Xpfet$151_0 vdd m1_31535_19792# vdd m1_17939_22513# pfet$151
Xnfet$179_3 m1_n10796_25662# m1_n9952_24224# m1_n8848_25658# vss nfet$179
Xnfet$158_8 m1_32193_25858# vss m1_32330_25662# vss nfet$158
Xpfet$142_27 vdd m1_14422_22513# m1_14422_22513# m1_14022_22402# m1_14556_21786# m1_14556_21786#
+ pfet$142
Xpfet$142_16 vdd m1_24973_22513# m1_24973_22513# m1_23945_22102# m1_25739_21786# m1_25739_21786#
+ pfet$142
Xnfet$184_1 m1_n5227_20152# vss m1_n6380_21786# vss nfet$184
Xnfet$177_0 m1_n8625_26174# vss m1_n8055_24542# vss nfet$177
Xpfet$169_1 vdd vdd vdd m1_n5019_22344# m1_n4485_21904# m1_n4485_21904# pfet$169
Xnfet$163_6 m1_354_22513# m1_354_22513# m1_31535_22102# m1_31535_22102# m1_31771_21430#
+ vss nfet$163
Xnfet$170_7 m1_n7401_15478# m1_n7401_15478# m1_n927_19404# m1_n927_19404# m1_n695_20470#
+ vss nfet$170
Xnfet$149_4 m1_12259_24224# m1_12259_24224# m1_11903_24542# m1_11903_24542# m1_12357_24542#
+ vss nfet$149
Xpfet$148_6 vdd vdd m1_n290_24224# m1_n910_23922# pfet$148
Xnfet$161_3 m1_326_24346# m1_326_24346# vss vss m1_n192_24542# vss nfet$161
Xnfet$154_2 m1_12805_21786# vss m1_12935_21590# vss nfet$154
Xpfet$146_3 vdd vdd m1_5901_19550# m1_649_17714# pfet$146
Xnfet$152_10 m1_9015_17714# m1_9015_17714# vss vss m1_14005_20470# vss nfet$152
Xpfet$140_93 vdd m1_28991_24224# m1_30095_25658# m1_28010_25858# pfet$140
Xpfet$140_82 vdd vdd m1_21241_24346# m1_n7513_20152# pfet$140
Xpfet$140_71 vdd vdd m1_11039_21786# m1_11760_25858# pfet$140
Xpfet$140_60 vdd vdd m1_20126_25858# m1_21241_24346# pfet$140
Xpfet$151_1 vdd vdd m1_30256_19792# m1_21456_22513# pfet$151
Xpfet$144_0 vdd vdd m1_n1133_21590# m1_n1263_21786# pfet$144
Xnfet$179_4 m1_n4623_25487# m1_n2567_23922# m1_n3184_24224# vss nfet$179
Xnfet$158_9 m1_n7513_20152# vss m1_33790_24346# vss nfet$158
Xpfet$142_28 vdd m1_14422_22513# m1_14422_22513# m1_13394_22102# m1_15188_21786# m1_15188_21786#
+ pfet$142
Xpfet$142_17 vdd m1_21456_22513# m1_21456_22513# m1_21056_22402# m1_21590_21786# m1_21590_21786#
+ pfet$142
Xnfet$177_1 m1_n8625_26174# vss m1_n7082_23622# vss nfet$177
Xpfet$169_2 vdd m1_n5764_21786# m1_n5764_21786# m1_n5019_22344# m1_n5227_21418# m1_n5227_21418#
+ pfet$169
Xnfet$163_7 m1_3871_22513# m1_3871_22513# vss vss m1_31771_21430# vss nfet$163
Xnfet$155_10 m1_26063_15478# vss m1_29239_20152# vss nfet$155
Xnfet$170_8 m1_26063_15478# m1_26063_15478# m1_n3822_20130# m1_n3822_20130# m1_27441_20470#
+ vss nfet$170
Xnfet$149_5 m1_8692_24346# m1_8692_24346# vss vss m1_8174_24542# vss nfet$149
Xpfet$148_7 vdd vdd m1_32330_25662# m1_32193_25858# pfet$148
Xnfet$161_4 m1_33174_24224# m1_33174_24224# m1_32818_24542# m1_32818_24542# m1_33272_24542#
+ vss nfet$161
Xpfet$146_4 vdd vdd m1_12935_19550# m1_9015_17714# pfet$146
Xnfet$154_3 m1_9288_21786# vss m1_9418_21590# vss nfet$154
Xnfet$152_11 m1_13198_17714# m1_13198_17714# vss vss m1_17522_20470# vss nfet$152
Xnfet$152_0 m1_n3534_17714# m1_n3534_17714# vss vss m1_3454_20470# vss nfet$152
Xpfet$151_2 vdd m1_30256_19792# vdd m1_24973_22513# pfet$151
Xpfet$144_1 vdd vdd m1_11671_21786# m1_11039_21786# pfet$144
Xpfet$140_94 vdd m1_28492_25858# vdd m1_30095_25658# pfet$140
Xpfet$140_83 vdd m1_21729_25658# m1_22522_24542# m1_19781_25662# pfet$140
Xpfet$140_72 vdd m1_13363_25658# m1_14156_24542# m1_11415_25662# pfet$140
Xpfet$140_61 vdd m1_24452_24542# vdd m1_25424_24346# pfet$140
Xpfet$140_50 vdd vdd m1_20268_25662# m1_20126_25858# pfet$140
Xnfet$158_10 m1_32675_25947# vss m1_35071_24542# vss nfet$158
Xnfet$179_5 m1_n4464_25980# m1_n3541_23922# m1_n4362_24346# vss nfet$179
Xnfet$169_20 m1_22493_16080# m1_22493_16080# m1_22034_17714# m1_22034_17714# m1_22591_16398#
+ vss nfet$169
Xnfet$177_2 vss vss m1_n9336_24346# vss nfet$177
Xpfet$142_29 vdd vdd vdd m1_14022_22402# m1_12805_21786# m1_12805_21786# pfet$142
Xpfet$142_18 vdd vdd vdd m1_24573_22402# m1_23356_21786# m1_23356_21786# pfet$142
Xnfet$155_11 m1_9331_15478# vss m1_15171_20152# vss nfet$155
Xnfet$170_9 m1_29239_20152# m1_29239_20152# m1_n3822_20130# m1_n3822_20130# m1_28073_20470#
+ vss nfet$170
Xnfet$149_6 m1_8076_24224# m1_8076_24224# m1_7720_24542# m1_7720_24542# m1_8174_24542#
+ vss nfet$149
Xpfet$148_8 vdd vdd m1_33174_24224# m1_32554_23922# pfet$148
Xnfet$182_0 m1_n4485_21904# m1_n5764_21786# vss vss nfet$182
Xpfet$167_0 vdd vdd m1_n7186_25858# m1_n10452_25858# pfet$167
Xnfet$161_5 m1_33790_24346# m1_33790_24346# vss vss m1_33272_24542# vss nfet$161
Xnfet$154_4 m1_7522_21786# vss m1_8154_21786# vss nfet$154
Xpfet$146_5 vdd vdd m1_8137_20152# m1_965_15478# pfet$146
Xnfet$152_12 m1_16452_19550# m1_16452_19550# vss vss m1_16890_20470# vss nfet$152
Xpfet$151_3 vdd vdd m1_34843_21786# m1_34093_19792# pfet$151
Xnfet$152_1 m1_2384_19550# m1_2384_19550# vss vss m1_2822_20470# vss nfet$152
Xpfet$144_2 vdd vdd m1_12935_21590# m1_12805_21786# pfet$144
Xpfet$140_95 vdd vdd m1_28991_24224# m1_28371_23922# pfet$140
Xpfet$140_84 vdd vdd m1_23827_25858# m1_18073_21786# pfet$140
Xpfet$140_73 vdd m1_16086_24542# vdd m1_17058_24346# pfet$140
Xpfet$140_62 vdd vdd m1_24452_24542# m1_24808_24224# pfet$140
Xpfet$140_51 vdd vdd m1_20625_24224# m1_20005_23922# pfet$140
Xpfet$140_40 vdd vdd m1_11760_25858# m1_12875_24346# pfet$140
Xnfet$158_11 m1_32554_23922# vss m1_33174_24224# vss nfet$158
Xnfet$179_6 m1_n4464_25980# m1_n3184_24224# m1_n3651_26174# vss nfet$179
Xnfet$169_10 m1_1578_16080# m1_1578_16080# m1_1119_17714# m1_1119_17714# m1_1676_16398#
+ vss nfet$169
Xnfet$177_3 fin vss m1_n10933_25858# vss nfet$177
Xpfet$142_19 vdd m1_24973_22513# m1_24973_22513# m1_24573_22402# m1_25107_21786# m1_25107_21786#
+ pfet$142
Xnfet$169_21 m1_14127_16080# m1_14127_16080# vss vss m1_15690_17358# vss nfet$169
Xnfet$149_7 m1_9180_25658# m1_9180_25658# vss vss m1_9639_25502# vss nfet$149
Xpfet$148_9 vdd vdd m1_28624_21786# m1_32675_25947# pfet$148
Xnfet$155_12 m1_13514_15478# vss m1_18688_20152# vss nfet$155
Xnfet$182_1 m1_n5227_21418# vss m1_n5764_21786# vss nfet$182
Xnfet$175_0 m1_n7082_23622# m1_n6856_24542# vss vss nfet$175
Xpfet$167_1 vdd m1_n7186_25858# vdd m1_n6111_25858# pfet$167
Xnfet$161_6 m1_33790_24346# m1_33790_24346# m1_32675_25947# m1_32675_25947# m1_34737_25502#
+ vss nfet$161
Xnfet$154_5 m1_488_21786# vss m1_1120_21786# vss nfet$154
Xpfet$146_6 vdd vdd m1_9418_19550# m1_4832_17714# pfet$146
Xnfet$152_13 m1_19969_19550# m1_19969_19550# vss vss m1_20407_20470# vss nfet$152
Xpfet$151_4 vdd m1_34093_19792# vdd m1_32818_20470# pfet$151
Xnfet$152_2 m1_5901_19550# m1_5901_19550# vss vss m1_6339_20470# vss nfet$152
Xnfet$177_10 vss vss m1_n4978_24224# vss nfet$177
Xpfet$144_3 vdd vdd m1_9418_21590# m1_9288_21786# pfet$144
Xpfet$140_96 vdd m1_28635_24542# vdd m1_29607_24346# pfet$140
Xpfet$140_85 vdd m1_24188_23922# m1_24452_24542# m1_23827_25858# pfet$140
Xpfet$140_74 vdd vdd m1_14556_21786# m1_15943_25858# pfet$140
Xpfet$140_63 vdd vdd m1_19781_25662# m1_19644_25858# pfet$140
Xpfet$140_52 vdd m1_20268_25662# m1_20005_23922# m1_19781_25662# pfet$140
Xpfet$140_41 vdd vdd m1_9288_21786# pd4 pfet$140
Xpfet$140_30 vdd vdd m1_2912_25858# m1_488_21786# pfet$140
Xpfet$142_0 vdd vdd vdd m1_n674_22102# m1_n1133_21590# m1_n1133_21590# pfet$142
Xnfet$158_12 m1_32675_25947# vss m1_28624_21786# vss nfet$158
Xnfet$179_7 m1_n4623_25487# m1_n4362_24346# m1_n4847_25662# vss nfet$179
Xpfet$141_110 vdd vdd m1_10458_17836# m1_10299_17343# pfet$141
Xnfet$169_22 m1_15564_15778# m1_15564_15778# m1_15454_18030# m1_15454_18030# m1_15690_17358#
+ vss nfet$169
Xnfet$169_11 m1_6377_16202# m1_6377_16202# vss vss m1_5859_16398# vss nfet$169
Xnfet$177_4 m1_n10572_23922# vss m1_n9952_24224# vss nfet$177
Xnfet$168_0 fout vss m1_35837_22102# vss nfet$168
Xnfet$155_13 m1_13198_17714# vss m1_16452_19550# vss nfet$155
Xnfet$149_8 m1_8692_24346# m1_8692_24346# m1_7577_25858# m1_7577_25858# m1_9639_25502#
+ vss nfet$149
Xnfet$182_2 m1_n6839_21786# vss m1_n6973_21481# vss nfet$182
Xnfet$175_1 m1_n8283_19850# vss m1_n6856_24542# vss nfet$175
Xpfet$143_30 vdd vdd vdd m1_24560_19550# m1_21880_15478# m1_21880_15478# pfet$143
Xnfet$161_7 m1_34278_25658# m1_34278_25658# vss vss m1_34737_25502# vss nfet$161
Xnfet$154_6 m1_5771_21786# vss m1_5901_21590# vss nfet$154
Xpfet$146_7 vdd vdd m1_11654_20152# m1_5148_15478# pfet$146
Xnfet$152_14 m1_17381_17714# m1_17381_17714# vss vss m1_21039_20470# vss nfet$152
Xpfet$172_0 vdd vdd m1_n8145_21908# m1_n6839_20152# pfet$172
Xnfet$152_3 m1_4832_17714# m1_4832_17714# vss vss m1_10488_20470# vss nfet$152
Xnfet$177_11 m1_n10452_25858# vss m1_n4847_25662# vss nfet$177
Xpfet$140_97 vdd vdd m1_21590_21786# m1_24309_25858# pfet$140
Xpfet$140_86 vdd m1_28634_25662# m1_28371_23922# m1_28147_25662# pfet$140
Xpfet$140_75 vdd vdd m1_19644_25858# m1_14556_21786# pfet$140
Xpfet$140_64 vdd vdd m1_22522_24542# m1_20126_25858# pfet$140
Xpfet$140_53 vdd m1_20625_24224# m1_21729_25658# m1_19644_25858# pfet$140
Xpfet$140_42 vdd m1_11760_25858# vdd m1_13363_25658# pfet$140
Xpfet$151_5 vdd vdd m1_34093_19792# m1_32818_21586# pfet$151
Xpfet$140_31 vdd m1_3273_23922# m1_3537_24542# m1_2912_25858# pfet$140
Xpfet$140_20 vdd vdd m1_4509_24346# m1_n7513_20152# pfet$140
Xpfet$144_4 vdd vdd m1_8154_21786# m1_7522_21786# pfet$144
Xpfet$142_1 vdd m1_7388_22513# m1_7388_22513# m1_6988_22402# m1_7522_21786# m1_7522_21786#
+ pfet$142
Xnfet$150_0 m1_3394_25858# vss m1_5790_24542# vss nfet$150
Xnfet$158_13 m1_32675_25947# vss m1_32817_25662# vss nfet$158
Xpfet$141_100 vdd vdd m1_23820_18030# m1_23930_15778# pfet$141
Xnfet$169_23 m1_18926_16202# m1_18926_16202# vss vss m1_18408_16398# vss nfet$169
Xnfet$169_12 m1_n1168_15778# m1_n1168_15778# m1_n1278_18030# m1_n1278_18030# m1_n1042_17358#
+ vss nfet$169
Xnfet$177_5 m1_n10933_25858# vss m1_n10796_25662# vss nfet$177
Xnfet$150_80 m1_28147_25662# m1_28991_24224# m1_30095_25658# vss nfet$150
Xnfet$149_9 m1_17058_24346# m1_17058_24346# vss vss m1_16540_24542# vss nfet$149
Xnfet$155_14 m1_21564_17714# vss m1_23486_19550# vss nfet$155
Xnfet$168_1 define m1_35837_22102# vss vss nfet$168
Xpfet$143_31 vdd m1_n2543_20130# m1_n2543_20130# m1_20407_19850# m1_19969_19550# m1_19969_19550#
+ pfet$143
Xpfet$143_20 vdd m1_n3822_21786# m1_n3822_21786# m1_14009_19550# m1_9015_17714# m1_9015_17714#
+ pfet$143
Xnfet$154_7 m1_4005_21786# vss m1_4637_21786# vss nfet$154
Xpfet$146_8 vdd vdd m1_n1133_19550# m1_n7383_17599# pfet$146
Xnfet$180_0 m1_n7186_25858# vss m1_n7320_25516# vss nfet$180
Xpfet$165_0 vdd vdd m1_n4485_20152# m1_n3822_20130# pfet$165
Xnfet$152_15 m1_21564_17714# m1_21564_17714# vss vss m1_24556_20470# vss nfet$152
Xnfet$152_4 m1_9418_19550# m1_9418_19550# vss vss m1_9856_20470# vss nfet$152
Xnfet$177_12 m1_n10452_25858# vss m1_n5571_25662# vss nfet$177
Xpfet$140_98 vdd m1_30095_25658# m1_30888_24542# m1_28147_25662# pfet$140
Xpfet$140_87 vdd vdd m1_28147_25662# m1_28010_25858# pfet$140
Xpfet$140_76 vdd m1_20005_23922# m1_20269_24542# m1_19644_25858# pfet$140
Xpfet$140_65 vdd vdd m1_18073_21786# m1_20126_25858# pfet$140
Xpfet$140_54 vdd vdd m1_24808_24224# m1_24188_23922# pfet$140
Xpfet$140_43 vdd vdd m1_12805_21786# pd5 pfet$140
Xpfet$151_6 vdd vdd m1_31535_19792# m1_14422_22513# pfet$151
Xpfet$140_32 vdd vdd m1_7720_24542# m1_8076_24224# pfet$140
Xpfet$140_21 vdd m1_7456_23922# m1_7720_24542# m1_7095_25858# pfet$140
Xpfet$140_10 vdd m1_8076_24224# m1_9180_25658# m1_7095_25858# pfet$140
Xpfet$144_5 vdd vdd m1_1120_21786# m1_488_21786# pfet$144
Xnfet$153_80 m1_18824_17836# m1_19747_15778# m1_18926_16202# vss nfet$153
Xpfet$142_2 vdd m1_7388_22513# m1_7388_22513# m1_6360_22102# m1_8154_21786# m1_8154_21786#
+ pfet$142
Xnfet$150_1 m1_2912_25858# m1_4997_25658# m1_5790_24542# vss nfet$150
Xpfet$141_101 vdd vdd m1_19637_18030# m1_19747_15778# pfet$141
Xnfet$169_24 m1_18310_16080# m1_18310_16080# m1_17851_17714# m1_17851_17714# m1_18408_16398#
+ vss nfet$169
Xnfet$169_13 m1_n2605_16080# m1_n2605_16080# vss vss m1_n1042_17358# vss nfet$169
Xnfet$177_6 m1_n10452_25858# vss m1_n10309_25662# vss nfet$177
Xnfet$150_81 m1_n7513_20152# vss m1_25424_24346# vss nfet$150
Xnfet$150_70 m1_21590_21786# vss m1_28010_25858# vss nfet$150
Xnfet$155_15 m1_17697_15478# vss m1_22205_20152# vss nfet$155
Xpfet$143_32 vdd m1_n2543_20130# m1_n2543_20130# m1_21043_19550# m1_17381_17714# m1_17381_17714#
+ pfet$143
Xpfet$143_21 vdd vdd vdd m1_13373_19850# m1_15171_20152# m1_15171_20152# pfet$143
Xpfet$143_10 vdd vdd vdd m1_9856_19850# m1_11654_20152# m1_11654_20152# pfet$143
Xpfet$146_9 vdd vdd m1_27003_19550# m1_25747_17714# pfet$146
Xnfet$173_0 m1_n5351_15778# m1_n5351_15778# m1_n5461_18030# m1_n5461_18030# m1_n5225_17358#
+ vss nfet$173
Xnfet$180_1 m1_n6856_24542# vss m1_n6111_25858# vss nfet$180
Xnfet$154_8 m1_2254_21786# vss m1_2384_21590# vss nfet$154
Xpfet$158_0 vdd vdd m1_n7247_17714# m1_n6788_16080# pfet$158
Xpfet$165_1 vdd m1_n4485_21904# vdd m1_9624_19404# pfet$165
Xnfet$152_16 m1_23486_19550# m1_23486_19550# vss vss m1_23924_20470# vss nfet$152
Xnfet$152_5 m1_649_17714# m1_649_17714# vss vss m1_6971_20470# vss nfet$152
Xnfet$177_13 fin vss m1_n4623_25487# vss nfet$177
Xpfet$151_7 vdd vdd m1_31535_22102# m1_354_22513# pfet$151
Xpfet$140_33 vdd vdd m1_7522_21786# m1_7577_25858# pfet$140
Xpfet$140_22 vdd vdd m1_3537_24542# m1_3893_24224# pfet$140
Xpfet$140_11 vdd vdd m1_7719_25662# m1_7577_25858# pfet$140
Xpfet$144_6 vdd vdd m1_5901_21590# m1_5771_21786# pfet$144
Xpfet$140_99 vdd vdd m1_26705_24542# m1_24309_25858# pfet$140
Xpfet$140_88 vdd vdd m1_28634_25662# m1_28492_25858# pfet$140
Xpfet$140_77 vdd vdd m1_20269_24542# m1_20625_24224# pfet$140
Xpfet$140_66 vdd vdd m1_15461_25858# m1_11039_21786# pfet$140
Xpfet$140_55 vdd m1_24451_25662# m1_24188_23922# m1_23964_25662# pfet$140
Xpfet$140_44 vdd m1_15943_25858# vdd m1_17546_25658# pfet$140
Xnfet$153_81 m1_13198_17714# vss m1_10299_17343# vss nfet$153
Xnfet$153_70 m1_n7513_20152# vss m1_18310_16080# vss nfet$153
Xnfet$150_2 m1_n7513_20152# vss m1_4509_24346# vss nfet$150
Xpfet$142_3 vdd m1_9645_21447# m1_9645_21447# m1_10505_22402# m1_11039_21786# m1_11039_21786#
+ pfet$142
Xpfet$146_10 vdd vdd m1_29239_20152# m1_26063_15478# pfet$146
Xpfet$140_0 vdd vdd m1_3049_25662# m1_2912_25858# pfet$140
Xpfet$141_102 vdd vdd m1_13198_17714# m1_13668_17714# pfet$141
Xnfet$169_25 m1_14743_16202# m1_14743_16202# vss vss m1_14225_16398# vss nfet$169
Xnfet$169_14 m1_n2605_16080# m1_n2605_16080# m1_n3064_17714# m1_n3064_17714# m1_n2507_16398#
+ vss nfet$169
Xnfet$177_7 m1_n7320_25516# vss m1_n2567_23922# vss nfet$177
Xnfet$150_82 m1_11415_25662# m1_12259_24224# m1_13363_25658# vss nfet$150
Xnfet$150_71 m1_28147_25662# m1_28371_23922# m1_28635_24542# vss nfet$150
Xnfet$150_60 pd6 vss m1_16322_21786# vss nfet$150
Xnfet$155_16 m1_17381_17714# vss m1_19969_19550# vss nfet$155
Xpfet$143_33 vdd m1_n3206_20274# m1_n3206_20274# m1_24560_19550# m1_21564_17714# m1_21564_17714#
+ pfet$143
Xpfet$143_22 vdd vdd vdd m1_14009_19550# m1_9331_15478# m1_9331_15478# pfet$143
Xpfet$143_11 vdd vdd vdd m1_10492_19550# m1_5148_15478# m1_5148_15478# pfet$143
Xnfet$154_9 m1_23356_21786# vss m1_23486_21590# vss nfet$154
Xnfet$166_0 m1_34093_19792# vss m1_34843_21786# vss nfet$166
Xnfet$173_1 m1_n6788_16080# m1_n6788_16080# vss vss m1_n5225_17358# vss nfet$173
Xpfet$158_1 vdd m1_n7247_17714# vdd m1_n6172_16202# pfet$158
Xpfet$165_2 vdd m1_n5227_21418# vdd m1_2590_19404# pfet$165
Xnfet$152_17 m1_12935_19550# m1_12935_19550# vss vss m1_13373_20470# vss nfet$152
Xnfet$152_6 m1_n1133_19550# m1_n1133_19550# vss vss m1_n695_20470# vss nfet$152
Xpfet$144_7 vdd vdd m1_4637_21786# m1_4005_21786# pfet$144
Xpfet$140_89 vdd vdd m1_19839_21786# pd7 pfet$140
Xpfet$140_78 vdd m1_20269_24542# vdd m1_21241_24346# pfet$140
Xpfet$140_67 vdd m1_15822_23922# m1_16086_24542# m1_15461_25858# pfet$140
Xpfet$140_56 vdd m1_24808_24224# m1_25912_25658# m1_23827_25858# pfet$140
Xpfet$140_45 vdd vdd m1_16442_24224# m1_15822_23922# pfet$140
Xpfet$140_34 vdd m1_9180_25658# m1_9973_24542# m1_7232_25662# pfet$140
Xpfet$140_23 vdd m1_3537_24542# vdd m1_4509_24346# pfet$140
Xpfet$140_12 vdd m1_7577_25858# vdd m1_9180_25658# pfet$140
Xpfet$170_0 vdd vdd m1_n5227_20152# m1_n2543_20130# pfet$170
Xnfet$150_3 m1_488_21786# vss m1_2912_25858# vss nfet$150
Xnfet$153_82 m1_10299_17343# vss m1_10458_17836# vss nfet$153
Xnfet$153_71 m1_14641_17836# m1_15921_16080# m1_15454_18030# vss nfet$153
Xnfet$153_60 m1_18665_17343# vss m1_18824_17836# vss nfet$153
Xpfet$142_4 vdd vdd vdd m1_9877_22102# m1_9418_21590# m1_9418_21590# pfet$142
Xpfet$141_103 vdd m1_14743_16202# m1_14258_17518# m1_14641_17836# pfet$141
Xpfet$146_11 vdd vdd m1_18688_20152# m1_13514_15478# pfet$146
Xnfet$169_26 m1_14127_16080# m1_14127_16080# m1_13668_17714# m1_13668_17714# m1_14225_16398#
+ vss nfet$169
Xpfet$140_1 vdd m1_3536_25662# m1_3273_23922# m1_3049_25662# pfet$140
Xnfet$169_15 m1_n1989_16202# m1_n1989_16202# vss vss m1_n2507_16398# vss nfet$169
Xnfet$177_8 m1_n4623_25487# vss m1_n4464_25980# vss nfet$177
Xnfet$150_72 m1_23827_25858# m1_25912_25658# m1_26705_24542# vss nfet$150
Xnfet$150_61 m1_23964_25662# m1_24808_24224# m1_25912_25658# vss nfet$150
Xnfet$150_50 m1_n7513_20152# vss m1_21241_24346# vss nfet$150
Xnfet$155_17 m1_21880_15478# vss m1_25722_20152# vss nfet$155
Xpfet$143_34 vdd m1_n3206_20274# m1_n3206_20274# m1_23924_19850# m1_23486_19550# m1_23486_19550#
+ pfet$143
Xpfet$143_23 vdd vdd vdd m1_16890_19850# m1_18688_20152# m1_18688_20152# pfet$143
Xpfet$143_12 vdd m1_6107_19404# m1_6107_19404# m1_6975_19550# m1_649_17714# m1_649_17714#
+ pfet$143
Xnfet$166_1 m1_30256_19792# vss m1_32818_20470# vss nfet$166
Xnfet$173_2 m1_n6788_16080# m1_n6788_16080# m1_n7247_17714# m1_n7247_17714# m1_n6690_16398#
+ vss nfet$173
Xpfet$165_3 vdd vdd m1_n5227_21418# m1_6107_19404# pfet$165
Xnfet$159_0 m1_n1134_25662# m1_n910_23922# m1_n646_24542# vss nfet$159
Xpfet$158_2 vdd vdd m1_n5461_18030# m1_n5351_15778# pfet$158
Xnfet$152_7 m1_n7383_17599# m1_n7383_17599# vss vss m1_n63_20470# vss nfet$152
Xpfet$144_8 vdd vdd m1_2384_21590# m1_2254_21786# pfet$144
Xpfet$140_79 vdd m1_17546_25658# m1_18339_24542# m1_15598_25662# pfet$140
Xpfet$140_68 vdd vdd m1_16086_24542# m1_16442_24224# pfet$140
Xpfet$140_57 vdd vdd m1_24451_25662# m1_24309_25858# pfet$140
Xpfet$140_46 vdd m1_16442_24224# m1_17546_25658# m1_15461_25858# pfet$140
Xpfet$140_35 vdd m1_7720_24542# vdd m1_8692_24346# pfet$140
Xpfet$140_24 vdd vdd m1_5790_24542# m1_3394_25858# pfet$140
Xpfet$140_13 vdd vdd m1_12259_24224# m1_11639_23922# pfet$140
Xpfet$170_1 vdd m1_n4485_20152# vdd m1_n3206_20274# pfet$170
Xpfet$163_0 vdd vdd m1_n7320_25516# m1_n7186_25858# pfet$163
Xnfet$150_4 m1_2912_25858# vss m1_3049_25662# vss nfet$150
Xnfet$153_72 m1_17851_17714# vss m1_18441_17518# vss nfet$153
Xnfet$153_61 m1_20104_16080# vss m1_19747_15778# vss nfet$153
Xnfet$153_50 m1_25747_17714# vss m1_22848_17343# vss nfet$153
Xpfet$142_5 vdd m1_9645_21447# m1_9645_21447# m1_9877_22102# m1_11671_21786# m1_11671_21786#
+ pfet$142
Xpfet$141_104 vdd vdd m1_14127_16080# m1_n7513_20152# pfet$141
Xpfet$146_12 vdd vdd m1_15171_20152# m1_9331_15478# pfet$146
Xpfet$140_2 vdd vdd m1_3394_25858# m1_4509_24346# pfet$140
Xnfet$150_62 m1_24188_23922# vss m1_24808_24224# vss nfet$150
Xnfet$150_51 m1_19644_25858# m1_21729_25658# m1_22522_24542# vss nfet$150
Xnfet$150_40 m1_15598_25662# m1_16442_24224# m1_17546_25658# vss nfet$150
Xnfet$169_27 m1_18310_16080# m1_18310_16080# vss vss m1_19873_17358# vss nfet$169
Xnfet$169_16 m1_19747_15778# m1_19747_15778# m1_19637_18030# m1_19637_18030# m1_19873_17358#
+ vss nfet$169
Xnfet$177_9 m1_n3184_24224# vss m1_n3541_23922# vss nfet$177
Xnfet$150_73 m1_24309_25858# vss m1_21590_21786# vss nfet$150
Xpfet$143_35 vdd m1_n3822_21786# m1_n3822_21786# m1_13373_19850# m1_12935_19550# m1_12935_19550#
+ pfet$143
Xpfet$143_24 vdd m1_n1927_20274# m1_n1927_20274# m1_16890_19850# m1_16452_19550# m1_16452_19550#
+ pfet$143
Xpfet$143_13 vdd m1_n927_19404# m1_n927_19404# m1_n695_19850# m1_n1133_19550# m1_n1133_19550#
+ pfet$143
Xnfet$166_2 m1_31535_19792# m1_32818_20470# vss vss nfet$166
Xnfet$173_3 m1_n6172_16202# m1_n6172_16202# vss vss m1_n6690_16398# vss nfet$173
Xnfet$159_1 m1_n1271_25858# m1_n647_25662# m1_n910_23922# vss nfet$159
Xpfet$158_3 vdd m1_n5461_18030# vdd m1_n6788_16080# pfet$158
Xpfet$165_4 vdd vdd m1_n4485_21904# m1_n3822_21786# pfet$165
Xnfet$152_8 m1_27003_19550# m1_27003_19550# vss vss m1_27441_20470# vss nfet$152
Xpfet$156_0 vdd vdd fout m1_34093_22102# pfet$156
Xpfet$140_69 vdd vdd m1_12875_24346# m1_n7513_20152# pfet$140
Xpfet$140_58 vdd vdd m1_23964_25662# m1_23827_25858# pfet$140
Xpfet$140_47 vdd vdd m1_15943_25858# m1_17058_24346# pfet$140
Xpfet$144_9 vdd vdd m1_22222_21786# m1_21590_21786# pfet$144
Xnfet$171_0 m1_35837_22102# vss m1_n7513_20152# vss nfet$171
Xpfet$140_36 vdd vdd m1_8692_24346# m1_n7513_20152# pfet$140
Xpfet$140_25 vdd vdd m1_4005_21786# m1_3394_25858# pfet$140
Xpfet$140_14 vdd vdd m1_11902_25662# m1_11760_25858# pfet$140
Xpfet$170_2 vdd m1_n5227_20152# vdd m1_n1927_20274# pfet$170
Xpfet$163_1 vdd vdd m1_n6111_25858# m1_n6856_24542# pfet$163
Xnfet$153_73 m1_13668_17714# vss m1_16538_15778# vss nfet$153
Xnfet$153_62 m1_18665_17343# m1_20721_15778# m1_20104_16080# vss nfet$153
Xnfet$153_51 m1_n7513_20152# vss m1_22493_16080# vss nfet$153
Xnfet$150_5 m1_2912_25858# m1_3536_25662# m1_3273_23922# vss nfet$150
Xnfet$153_40 m1_n2250_17343# m1_n194_15778# m1_n811_16080# vss nfet$153
Xpfet$142_6 vdd vdd vdd m1_10505_22402# m1_9288_21786# m1_9288_21786# pfet$142
Xpfet$141_90 vdd m1_19747_15778# m1_18926_16202# m1_18665_17343# pfet$141
Xpfet$146_13 vdd vdd m1_16452_19550# m1_13198_17714# pfet$146
Xpfet$140_3 vdd m1_3394_25858# vdd m1_4997_25658# pfet$140
Xpfet$141_105 vdd vdd m1_14258_17518# m1_13668_17714# pfet$141
Xnfet$169_17 m1_22493_16080# m1_22493_16080# vss vss m1_24056_17358# vss nfet$169
Xnfet$150_74 pd8 vss m1_23356_21786# vss nfet$150
Xnfet$150_63 m1_14556_21786# vss m1_19644_25858# vss nfet$150
Xnfet$150_52 m1_20126_25858# vss m1_22522_24542# vss nfet$150
Xnfet$150_41 pd5 vss m1_12805_21786# vss nfet$150
Xnfet$150_30 m1_n7513_20152# vss m1_17058_24346# vss nfet$150
Xpfet$143_25 vdd vdd vdd m1_17526_19550# m1_13514_15478# m1_13514_15478# pfet$143
Xpfet$143_14 vdd m1_n927_19404# m1_n927_19404# m1_n59_19550# m1_n7383_17599# m1_n7383_17599#
+ pfet$143
Xnfet$166_3 m1_30256_22102# vss m1_32818_21586# vss nfet$166
Xnfet$173_4 m1_28113_15778# m1_28113_15778# m1_28003_18030# m1_28003_18030# m1_28239_17358#
+ vss nfet$173
Xnfet$159_2 m1_n1271_25858# m1_814_25658# m1_1607_24542# vss nfet$159
Xpfet$158_4 vdd vdd m1_26217_17714# m1_26676_16080# pfet$158
Xpfet$165_5 vdd m1_n6839_21786# vdd m1_n5764_21786# pfet$165
Xnfet$152_9 m1_25747_17714# m1_25747_17714# vss vss m1_28073_20470# vss nfet$152
Xnfet$164_0 m1_34843_21786# m1_34843_21786# m1_34093_22102# m1_34093_22102# m1_34329_21430#
+ vss nfet$164
Xpfet$140_59 vdd vdd m1_16322_21786# pd6 pfet$140
Xpfet$140_48 vdd m1_16085_25662# m1_15822_23922# m1_15598_25662# pfet$140
Xpfet$140_37 vdd vdd m1_9973_24542# m1_7577_25858# pfet$140
Xpfet$140_26 vdd m1_4997_25658# m1_5790_24542# m1_3049_25662# pfet$140
Xpfet$140_15 vdd m1_11902_25662# m1_11639_23922# m1_11415_25662# pfet$140
Xpfet$170_3 vdd m1_n6839_20152# vdd m1_n927_19404# pfet$170
Xpfet$149_0 vdd vdd m1_n646_24542# m1_n290_24224# pfet$149
Xnfet$153_74 m1_14482_17343# vss m1_14641_17836# vss nfet$153
Xnfet$153_63 m1_13668_17714# vss m1_14258_17518# vss nfet$153
Xnfet$153_52 m1_23007_17836# m1_24287_16080# m1_23820_18030# vss nfet$153
Xnfet$150_6 m1_3049_25662# m1_3893_24224# m1_4997_25658# vss nfet$150
Xnfet$153_30 sd6 vss m1_5148_15478# vss nfet$153
Xnfet$153_41 m1_n2091_17836# m1_n1168_15778# m1_n1989_16202# vss nfet$153
Xpfet$142_7 vdd m1_354_22513# m1_354_22513# m1_n674_22102# m1_1120_21786# m1_1120_21786#
+ pfet$142
Xpfet$141_91 vdd m1_24287_16080# m1_23820_18030# m1_22848_17343# pfet$141
Xpfet$141_80 vdd vdd m1_15564_15778# m1_15921_16080# pfet$141
Xpfet$146_14 vdd vdd m1_23486_19550# m1_21564_17714# pfet$146
Xpfet$140_4 vdd vdd m1_3893_24224# m1_3273_23922# pfet$140
Xpfet$141_106 vdd vdd m1_14482_17343# m1_17381_17714# pfet$141
Xnfet$169_18 m1_23930_15778# m1_23930_15778# m1_23820_18030# m1_23820_18030# m1_24056_17358#
+ vss nfet$169
Xnfet$150_75 m1_28371_23922# vss m1_28991_24224# vss nfet$150
Xnfet$150_64 m1_19644_25858# vss m1_19781_25662# vss nfet$150
Xnfet$150_53 m1_23827_25858# m1_24451_25662# m1_24188_23922# vss nfet$150
Xnfet$150_42 m1_15943_25858# vss m1_16085_25662# vss nfet$150
Xnfet$150_31 m1_15943_25858# vss m1_18339_24542# vss nfet$150
Xnfet$150_20 pd3 vss m1_5771_21786# vss nfet$150
Xpfet$143_26 vdd m1_n1927_20274# m1_n1927_20274# m1_17526_19550# m1_13198_17714# m1_13198_17714#
+ pfet$143
Xpfet$143_15 vdd vdd vdd m1_n59_19550# m1_n7401_15478# m1_n7401_15478# pfet$143
Xnfet$173_5 m1_26676_16080# m1_26676_16080# vss vss m1_28239_17358# vss nfet$173
Xpfet$158_5 vdd m1_26217_17714# vdd m1_27292_16202# pfet$158
Xnfet$159_3 m1_n1134_25662# m1_n290_24224# m1_814_25658# vss nfet$159
Xpfet$165_6 vdd vdd m1_n6973_21481# m1_n6839_21786# pfet$165
Xnfet$164_1 m1_28490_22513# m1_28490_22513# vss vss m1_34329_21430# vss nfet$164
Xpfet$140_49 vdd m1_20126_25858# vdd m1_21729_25658# pfet$140
Xpfet$140_38 vdd vdd m1_16085_25662# m1_15943_25858# pfet$140
Xpfet$140_27 vdd vdd m1_11278_25858# m1_7522_21786# pfet$140
Xpfet$140_16 vdd vdd m1_5771_21786# pd3 pfet$140
Xnfet$157_0 m1_n3534_17714# vss m1_n6433_17343# vss nfet$157
Xpfet$149_1 vdd m1_n789_25858# vdd m1_814_25658# pfet$149
Xpfet$170_4 vdd vdd m1_n6839_20152# m1_n6973_21481# pfet$170
Xnfet$153_75 sd3 vss m1_17697_15478# vss nfet$153
Xnfet$153_64 m1_13668_17714# vss m1_13198_17714# vss nfet$153
Xnfet$153_53 m1_22848_17343# vss m1_23007_17836# vss nfet$153
Xnfet$150_7 m1_3049_25662# m1_3273_23922# m1_3537_24542# vss nfet$150
Xnfet$153_31 m1_1933_17343# m1_3989_15778# m1_3372_16080# vss nfet$153
Xnfet$153_20 m1_1119_17714# vss m1_1709_17518# vss nfet$153
Xnfet$153_42 m1_n811_16080# vss m1_n1168_15778# vss nfet$153
Xpfet$161_0 vdd vdd vdd m1_n6624_23622# m1_n7082_23622# m1_n7082_23622# pfet$161
Xpfet$142_8 vdd vdd vdd m1_6360_22102# m1_5901_21590# m1_5901_21590# pfet$142
Xpfet$141_92 vdd m1_15454_18030# vdd m1_14127_16080# pfet$141
Xpfet$141_81 vdd vdd m1_13668_17714# m1_14127_16080# pfet$141
Xpfet$141_70 vdd vdd m1_18824_17836# m1_18665_17343# pfet$141
Xpfet$146_15 vdd vdd m1_22205_20152# m1_17697_15478# pfet$146
Xpfet$140_5 vdd m1_3893_24224# m1_4997_25658# m1_2912_25858# pfet$140
Xpfet$141_107 vdd m1_15921_16080# m1_15454_18030# m1_14482_17343# pfet$141
Xnfet$169_19 m1_23109_16202# m1_23109_16202# vss vss m1_22591_16398# vss nfet$169
Xnfet$150_76 m1_28492_25858# vss m1_28634_25662# vss nfet$150
Xnfet$150_65 m1_28492_25858# vss m1_25107_21786# vss nfet$150
Xnfet$150_54 m1_24309_25858# vss m1_24451_25662# vss nfet$150
Xnfet$150_43 m1_15461_25858# vss m1_15598_25662# vss nfet$150
Xnfet$150_32 m1_15461_25858# m1_17546_25658# m1_18339_24542# vss nfet$150
Xnfet$150_21 m1_11278_25858# m1_11902_25662# m1_11639_23922# vss nfet$150
Xnfet$150_10 m1_7577_25858# vss m1_9973_24542# vss nfet$150
Xpfet$143_27 vdd vdd vdd m1_20407_19850# m1_22205_20152# m1_22205_20152# pfet$143
Xpfet$143_16 vdd vdd vdd m1_28077_19550# m1_26063_15478# m1_26063_15478# pfet$143
Xnfet$159_4 m1_32193_25858# m1_34278_25658# m1_35071_24542# vss nfet$159
Xpfet$158_6 vdd vdd m1_28003_18030# m1_28113_15778# pfet$158
Xnfet$173_6 m1_27292_16202# m1_27292_16202# vss vss m1_26774_16398# vss nfet$173
Xpfet$165_7 vdd vdd m1_n6839_21786# m1_n6380_21786# pfet$165
Xnfet$164_2 m1_9645_21447# m1_9645_21447# vss vss m1_30492_21430# vss nfet$164
Xnfet$157_1 m1_n7513_20152# vss m1_n6788_16080# vss nfet$157
Xpfet$140_39 vdd vdd m1_15598_25662# m1_15461_25858# pfet$140
Xpfet$140_28 vdd m1_11639_23922# m1_11903_24542# m1_11278_25858# pfet$140
Xpfet$140_17 vdd vdd m1_7577_25858# m1_8692_24346# pfet$140
Xpfet$149_2 vdd vdd m1_n789_25858# m1_326_24346# pfet$149
Xnfet$150_8 m1_3394_25858# vss m1_3536_25662# vss nfet$150
Xnfet$153_76 m1_14482_17343# m1_16538_15778# m1_15921_16080# vss nfet$153
Xnfet$153_65 m1_14482_17343# m1_14743_16202# m1_14258_17518# vss nfet$153
Xnfet$153_54 m1_22848_17343# m1_23109_16202# m1_22624_17518# vss nfet$153
Xnfet$153_32 m1_2092_17836# m1_3015_15778# m1_2194_16202# vss nfet$153
Xnfet$153_21 m1_1933_17343# m1_2194_16202# m1_1709_17518# vss nfet$153
Xnfet$153_10 m1_11738_16080# vss m1_11381_15778# vss nfet$153
Xnfet$153_43 sd8 vss m1_n3218_15478# vss nfet$153
Xpfet$142_9 vdd m1_3871_22513# m1_3871_22513# m1_3471_22402# m1_4005_21786# m1_4005_21786#
+ pfet$142
Xpfet$154_0 vdd m1_34093_22102# vdd m1_28490_22513# pfet$154
Xpfet$141_93 vdd m1_23820_18030# vdd m1_22493_16080# pfet$141
Xpfet$141_82 vdd m1_13668_17714# vdd m1_14743_16202# pfet$141
Xpfet$141_71 vdd vdd m1_19747_15778# m1_20104_16080# pfet$141
Xpfet$141_60 vdd vdd m1_n194_15778# m1_n3064_17714# pfet$141
Xpfet$161_1 vdd m1_n6856_24542# m1_n6856_24542# m1_n6624_23622# m1_n8283_19850# m1_n8283_19850#
+ pfet$161
Xpfet$141_108 vdd vdd m1_15454_18030# m1_15564_15778# pfet$141
Xpfet$146_16 vdd vdd m1_19969_19550# m1_17381_17714# pfet$146
Xpfet$140_6 vdd vdd m1_3536_25662# m1_3394_25858# pfet$140
Xnfet$150_77 m1_28010_25858# vss m1_28147_25662# vss nfet$150
Xnfet$150_66 m1_28010_25858# m1_30095_25658# m1_30888_24542# vss nfet$150
Xnfet$150_55 m1_23827_25858# vss m1_23964_25662# vss nfet$150
Xnfet$150_44 m1_15822_23922# vss m1_16442_24224# vss nfet$150
Xnfet$150_33 m1_11760_25858# vss m1_14156_24542# vss nfet$150
Xnfet$150_22 m1_11760_25858# vss m1_11902_25662# vss nfet$150
Xnfet$150_11 m1_7522_21786# vss m1_11278_25858# vss nfet$150
Xpfet$143_28 vdd vdd vdd m1_21043_19550# m1_17697_15478# m1_17697_15478# pfet$143
Xpfet$143_17 vdd m1_n3822_20130# m1_n3822_20130# m1_28077_19550# m1_25747_17714# m1_25747_17714#
+ pfet$143
Xnfet$159_5 m1_32330_25662# m1_33174_24224# m1_34278_25658# vss nfet$159
Xnfet$173_7 m1_26676_16080# m1_26676_16080# m1_26217_17714# m1_26217_17714# m1_26774_16398#
+ vss nfet$173
Xpfet$158_7 vdd m1_28003_18030# vdd m1_26676_16080# pfet$158
Xnfet$164_3 m1_7388_22513# m1_7388_22513# m1_30256_22102# m1_30256_22102# m1_30492_21430#
+ vss nfet$164
Xpfet$149_3 vdd m1_n646_24542# vdd m1_326_24346# pfet$149
Xpfet$140_29 vdd vdd m1_11903_24542# m1_12259_24224# pfet$140
Xpfet$140_18 vdd vdd m1_11415_25662# m1_11278_25858# pfet$140
Xnfet$157_2 m1_n4994_16080# vss m1_n5351_15778# vss nfet$157
Xnfet$150_9 m1_3273_23922# vss m1_3893_24224# vss nfet$150
Xnfet$153_77 sd4 vss m1_13514_15478# vss nfet$153
Xnfet$153_66 m1_n7513_20152# vss m1_14127_16080# vss nfet$153
Xnfet$153_55 m1_22034_17714# vss m1_24904_15778# vss nfet$153
Xnfet$153_44 m1_n2091_17836# m1_n811_16080# m1_n1278_18030# vss nfet$153
Xnfet$153_33 sd7 vss m1_965_15478# vss nfet$153
Xnfet$153_22 m1_6116_17343# m1_6377_16202# m1_5892_17518# vss nfet$153
Xnfet$153_11 m1_10299_17343# m1_12355_15778# m1_11738_16080# vss nfet$153
Xnfet$162_0 m1_11039_21786# m1_11039_21786# vss vss m1_9877_21586# vss nfet$162
Xpfet$154_1 vdd vdd m1_34093_22102# m1_34843_21786# pfet$154
Xpfet$141_94 vdd vdd m1_22624_17518# m1_22034_17714# pfet$141
Xpfet$141_83 vdd m1_16538_15778# m1_15921_16080# m1_14641_17836# pfet$141
Xpfet$141_72 vdd m1_20721_15778# m1_20104_16080# m1_18824_17836# pfet$141
Xpfet$141_61 vdd m1_n811_16080# m1_n1278_18030# m1_n2250_17343# pfet$141
Xpfet$141_50 vdd m1_n1168_15778# m1_n1989_16202# m1_n2250_17343# pfet$141
Xpfet$147_0 vdd vdd m1_n7401_15478# sd9 pfet$147
Xpfet$141_109 vdd vdd m1_10299_17343# m1_13198_17714# pfet$141
Xpfet$146_17 vdd vdd m1_25722_20152# m1_21880_15478# pfet$146
Xpfet$140_7 vdd vdd m1_7232_25662# m1_7095_25858# pfet$140
Xnfet$150_78 m1_28010_25858# m1_28634_25662# m1_28371_23922# vss nfet$150
Xnfet$150_67 m1_28492_25858# vss m1_30888_24542# vss nfet$150
Xnfet$150_56 m1_19781_25662# m1_20625_24224# m1_21729_25658# vss nfet$150
Xnfet$150_45 m1_15461_25858# m1_16085_25662# m1_15822_23922# vss nfet$150
Xnfet$150_34 m1_11278_25858# m1_13363_25658# m1_14156_24542# vss nfet$150
Xnfet$150_23 m1_11278_25858# vss m1_11415_25662# vss nfet$150
Xnfet$150_12 m1_7577_25858# vss m1_7522_21786# vss nfet$150
Xpfet$143_29 vdd vdd vdd m1_23924_19850# m1_25722_20152# m1_25722_20152# pfet$143
Xpfet$143_18 vdd vdd vdd m1_27441_19850# m1_29239_20152# m1_29239_20152# pfet$143
Xnfet$159_6 m1_32193_25858# m1_32817_25662# m1_32554_23922# vss nfet$159
Xpfet$149_4 vdd vdd m1_32675_25947# m1_33790_24346# pfet$149
Xpfet$140_19 vdd vdd m1_7095_25858# m1_4005_21786# pfet$140
Xnfet$157_3 m1_n6433_17343# vss m1_n6274_17836# vss nfet$157
Xnfet$153_78 m1_14641_17836# m1_15564_15778# m1_14743_16202# vss nfet$153
Xnfet$153_67 m1_17381_17714# vss m1_14482_17343# vss nfet$153
Xnfet$153_56 m1_24287_16080# vss m1_23930_15778# vss nfet$153
Xnfet$153_45 m1_n3064_17714# vss m1_n194_15778# vss nfet$153
Xnfet$155_0 m1_n3534_17714# vss m1_2384_19550# vss nfet$155
Xnfet$153_34 m1_n2250_17343# vss m1_n2091_17836# vss nfet$153
Xnfet$153_23 m1_5302_17714# vss m1_4832_17714# vss nfet$153
Xnfet$153_12 m1_9485_17714# vss m1_12355_15778# vss nfet$153
Xnfet$162_1 m1_11671_21786# m1_11671_21786# vss vss m1_10509_21586# vss nfet$162
Xpfet$154_2 vdd vdd m1_30256_22102# m1_7388_22513# pfet$154
Xpfet$147_1 vdd vdd m1_21880_15478# sd2 pfet$147
Xpfet$141_95 vdd vdd m1_21564_17714# m1_22034_17714# pfet$141
Xpfet$141_84 vdd vdd m1_17381_17714# m1_17851_17714# pfet$141
Xpfet$141_73 vdd vdd m1_16538_15778# m1_13668_17714# pfet$141
Xpfet$141_62 vdd vdd m1_23007_17836# m1_22848_17343# pfet$141
Xpfet$141_40 vdd m1_10560_16202# m1_10075_17518# m1_10458_17836# pfet$141
Xpfet$141_51 vdd vdd m1_n1168_15778# m1_n811_16080# pfet$141
Xpfet$140_8 vdd vdd m1_8076_24224# m1_7456_23922# pfet$140
Xpfet$140_110 vdd m1_11903_24542# vdd m1_12875_24346# pfet$140
Xnfet$150_79 pd7 vss m1_19839_21786# vss nfet$150
Xnfet$150_68 m1_n7513_20152# vss m1_29607_24346# vss nfet$150
Xnfet$150_57 m1_20126_25858# vss m1_20268_25662# vss nfet$150
Xnfet$150_46 m1_20126_25858# vss m1_18073_21786# vss nfet$150
Xnfet$150_35 m1_15598_25662# m1_15822_23922# m1_16086_24542# vss nfet$150
Xnfet$150_24 m1_7095_25858# m1_7719_25662# m1_7456_23922# vss nfet$150
Xnfet$150_13 m1_11415_25662# m1_11639_23922# m1_11903_24542# vss nfet$150
Xpfet$143_19 vdd m1_n3822_20130# m1_n3822_20130# m1_27441_19850# m1_27003_19550# m1_27003_19550#
+ pfet$143
Xnfet$159_7 m1_32330_25662# m1_32554_23922# m1_32818_24542# vss nfet$159
Xnfet$185_0 m1_n6839_20152# vss m1_n8145_21908# vss nfet$185
Xnfet$157_4 m1_n7247_17714# vss m1_n4377_15778# vss nfet$157
Xpfet$149_5 vdd m1_32675_25947# vdd m1_34278_25658# pfet$149
Xnfet$153_79 m1_15921_16080# vss m1_15564_15778# vss nfet$153
Xnfet$153_68 m1_18665_17343# m1_18926_16202# m1_18441_17518# vss nfet$153
Xnfet$153_57 m1_22848_17343# m1_24904_15778# m1_24287_16080# vss nfet$153
Xnfet$153_46 m1_22034_17714# vss m1_21564_17714# vss nfet$153
Xnfet$153_24 m1_4832_17714# vss m1_1933_17343# vss nfet$153
Xnfet$153_13 m1_10458_17836# m1_11381_15778# m1_10560_16202# vss nfet$153
Xnfet$153_35 m1_n7513_20152# vss m1_5761_16080# vss nfet$153
Xpfet$147_2 vdd vdd m1_26063_15478# sd1 pfet$147
Xpfet$154_3 vdd m1_31535_22102# vdd m1_3871_22513# pfet$154
Xnfet$155_1 m1_n3218_15478# vss m1_4620_20152# vss nfet$155
Xnfet$162_2 m1_8154_21786# m1_8154_21786# vss vss m1_6992_21586# vss nfet$162
Xpfet$141_96 vdd vdd m1_18665_17343# m1_21564_17714# pfet$141
Xpfet$141_85 vdd m1_18926_16202# m1_18441_17518# m1_18824_17836# pfet$141
Xpfet$141_74 vdd vdd m1_14641_17836# m1_14482_17343# pfet$141
Xpfet$141_63 vdd m1_23930_15778# m1_23109_16202# m1_22848_17343# pfet$141
Xpfet$141_30 vdd vdd m1_1933_17343# m1_4832_17714# pfet$141
Xpfet$141_41 vdd vdd m1_10075_17518# m1_9485_17714# pfet$141
Xpfet$141_52 vdd m1_n3064_17714# vdd m1_n1989_16202# pfet$141
Xpfet$140_9 vdd m1_7719_25662# m1_7456_23922# m1_7232_25662# pfet$140
Xpfet$152_0 vdd m1_n647_25662# m1_n910_23922# m1_n1134_25662# pfet$152
Xpfet$140_100 vdd vdd m1_29607_24346# m1_n7513_20152# pfet$140
Xnfet$150_69 m1_24309_25858# vss m1_26705_24542# vss nfet$150
Xnfet$150_58 m1_20005_23922# vss m1_20625_24224# vss nfet$150
Xnfet$150_47 m1_23964_25662# m1_24188_23922# m1_24452_24542# vss nfet$150
Xnfet$150_36 m1_11760_25858# vss m1_11039_21786# vss nfet$150
Xnfet$150_25 m1_7232_25662# m1_8076_24224# m1_9180_25658# vss nfet$150
Xnfet$150_14 m1_n7513_20152# vss m1_8692_24346# vss nfet$150
Xnfet$178_0 m1_n9952_24224# m1_n9952_24224# m1_n10308_24542# m1_n10308_24542# m1_n9854_24542#
+ vss nfet$178
Xnfet$157_5 m1_n7247_17714# vss m1_n6657_17518# vss nfet$157
Xpfet$149_6 vdd vdd m1_32818_24542# m1_33174_24224# pfet$149
Xnfet$153_69 m1_17851_17714# vss m1_17381_17714# vss nfet$153
Xnfet$153_58 m1_23007_17836# m1_23930_15778# m1_23109_16202# vss nfet$153
Xnfet$153_47 m1_22034_17714# vss m1_22624_17518# vss nfet$153
Xnfet$153_25 m1_2092_17836# m1_3372_16080# m1_2905_18030# vss nfet$153
Xnfet$153_14 m1_6116_17343# m1_8172_15778# m1_7555_16080# vss nfet$153
Xnfet$153_36 m1_n3064_17714# vss m1_n2474_17518# vss nfet$153
Xpfet$154_4 vdd m1_30256_22102# vdd m1_9645_21447# pfet$154
Xnfet$155_2 m1_n7401_15478# vss m1_1103_20152# vss nfet$155
Xnfet$162_3 m1_7522_21786# m1_7522_21786# vss vss m1_6360_21586# vss nfet$162
Xpfet$141_97 vdd vdd m1_22493_16080# m1_n7513_20152# pfet$141
Xpfet$141_86 vdd m1_19637_18030# vdd m1_18310_16080# pfet$141
Xpfet$141_75 vdd vdd m1_17697_15478# sd3 pfet$141
Xpfet$141_64 vdd vdd m1_23930_15778# m1_24287_16080# pfet$141
Xpfet$141_20 vdd vdd m1_1119_17714# m1_1578_16080# pfet$141
Xpfet$141_31 vdd m1_3372_16080# m1_2905_18030# m1_1933_17343# pfet$141
Xpfet$141_42 vdd m1_11271_18030# vdd m1_9944_16080# pfet$141
Xpfet$141_53 vdd vdd m1_n3218_15478# sd8 pfet$141
Xnfet$160_0 pd1 vss m1_n1263_21786# vss nfet$160
Xpfet$145_0 vdd vdd m1_n6274_17836# m1_n6433_17343# pfet$145
Xpfet$152_1 vdd m1_n910_23922# m1_n646_24542# m1_n1271_25858# pfet$152
Xpfet$140_101 vdd vdd m1_28010_25858# m1_21590_21786# pfet$140
Xnfet$150_59 m1_19644_25858# m1_20268_25662# m1_20005_23922# vss nfet$150
Xnfet$150_48 m1_18073_21786# vss m1_23827_25858# vss nfet$150
Xnfet$150_37 m1_11039_21786# vss m1_15461_25858# vss nfet$150
Xnfet$150_26 m1_7095_25858# m1_9180_25658# m1_9973_24542# vss nfet$150
Xnfet$150_15 m1_7232_25662# m1_7456_23922# m1_7720_24542# vss nfet$150
Xnfet$178_1 m1_n9336_24346# m1_n9336_24346# m1_n8625_26174# m1_n8625_26174# m1_n8389_25502#
+ vss nfet$178
Xnfet$157_6 m1_n7247_17714# vss m1_n7383_17599# vss nfet$157
Xpfet$149_7 vdd m1_32818_24542# vdd m1_33790_24346# pfet$149
Xnfet$153_59 m1_17851_17714# vss m1_20721_15778# vss nfet$153
Xnfet$153_48 m1_18824_17836# m1_20104_16080# m1_19637_18030# vss nfet$153
Xnfet$155_3 m1_649_17714# vss m1_5901_19550# vss nfet$155
Xnfet$153_26 m1_5302_17714# vss m1_5892_17518# vss nfet$153
Xnfet$153_15 m1_5302_17714# vss m1_8172_15778# vss nfet$153
Xnfet$153_37 m1_n7513_20152# vss m1_n2605_16080# vss nfet$153
Xnfet$162_4 m1_1120_21786# m1_1120_21786# vss vss m1_n42_21586# vss nfet$162
Xpfet$141_98 vdd m1_20104_16080# m1_19637_18030# m1_18665_17343# pfet$141
Xpfet$141_87 vdd vdd m1_18310_16080# m1_n7513_20152# pfet$141
Xpfet$141_76 vdd m1_17851_17714# vdd m1_18926_16202# pfet$141
Xpfet$141_65 vdd m1_24904_15778# m1_24287_16080# m1_23007_17836# pfet$141
Xpfet$141_21 vdd vdd m1_965_15478# sd7 pfet$141
Xpfet$141_10 vdd m1_8172_15778# m1_7555_16080# m1_6275_17836# pfet$141
Xpfet$141_32 vdd vdd m1_2905_18030# m1_3015_15778# pfet$141
Xpfet$141_43 vdd vdd m1_11271_18030# m1_11381_15778# pfet$141
Xpfet$141_54 vdd vdd m1_n1278_18030# m1_n1168_15778# pfet$141
Xnfet$160_1 pd2 vss m1_2254_21786# vss nfet$160
Xnfet$153_0 m1_9485_17714# vss m1_9015_17714# vss nfet$153
Xpfet$145_1 vdd vdd m1_n4377_15778# m1_n7247_17714# pfet$145
Xpfet$152_2 vdd m1_n290_24224# m1_814_25658# m1_n1271_25858# pfet$152
Xpfet$140_102 vdd m1_28371_23922# m1_28635_24542# m1_28010_25858# pfet$140
Xnfet$150_49 m1_19781_25662# m1_20005_23922# m1_20269_24542# vss nfet$150
Xnfet$150_38 m1_n7513_20152# vss m1_12875_24346# vss nfet$150
Xnfet$150_27 m1_7577_25858# vss m1_7719_25662# vss nfet$150
Xnfet$150_16 m1_4005_21786# vss m1_7095_25858# vss nfet$150
Xnfet$178_2 m1_n8848_25658# m1_n8848_25658# vss vss m1_n8389_25502# vss nfet$178
Xpfet$144_10 vdd vdd m1_23486_21590# m1_23356_21786# pfet$144
Xnfet$157_7 m1_26217_17714# vss m1_26807_17518# vss nfet$157
Xnfet$183_0 m1_n927_19404# m1_n927_19404# vss vss m1_n6282_20470# vss nfet$183
Xpfet$168_0 vdd vdd vdd m1_n8047_19550# m1_n7513_20152# m1_n7513_20152# pfet$168
Xnfet$153_49 m1_21564_17714# vss m1_18665_17343# vss nfet$153
Xnfet$155_4 m1_4832_17714# vss m1_9418_19550# vss nfet$155
Xnfet$153_27 m1_1119_17714# vss m1_3989_15778# vss nfet$153
Xnfet$153_16 m1_6275_17836# m1_7198_15778# m1_6377_16202# vss nfet$153
Xnfet$153_38 m1_n2250_17343# m1_n1989_16202# m1_n2474_17518# vss nfet$153
Xnfet$162_5 m1_4005_21786# m1_4005_21786# vss vss m1_2843_21586# vss nfet$162
Xpfet$141_99 vdd m1_23109_16202# m1_22624_17518# m1_23007_17836# pfet$141
Xpfet$141_88 vdd vdd m1_18441_17518# m1_17851_17714# pfet$141
Xpfet$141_77 vdd vdd m1_17851_17714# m1_18310_16080# pfet$141
Xpfet$141_66 vdd vdd m1_24904_15778# m1_22034_17714# pfet$141
Xpfet$141_22 vdd vdd m1_3015_15778# m1_3372_16080# pfet$141
Xpfet$141_11 vdd vdd m1_9485_17714# m1_9944_16080# pfet$141
Xpfet$141_33 vdd vdd m1_5892_17518# m1_5302_17714# pfet$141
Xpfet$141_44 vdd vdd m1_649_17714# m1_1119_17714# pfet$141
Xpfet$141_55 vdd vdd m1_n2474_17518# m1_n3064_17714# pfet$141
Xnfet$160_2 pd9 vss m1_26873_21786# vss nfet$160
Xnfet$153_1 m1_9015_17714# vss m1_6116_17343# vss nfet$153
Xpfet$140_103 vdd vdd m1_28635_24542# m1_28991_24224# pfet$140
Xnfet$150_39 pd4 vss m1_9288_21786# vss nfet$150
Xpfet$152_3 vdd m1_814_25658# m1_1607_24542# m1_n1134_25662# pfet$152
Xnfet$150_28 m1_3394_25858# vss m1_4005_21786# vss nfet$150
Xnfet$150_17 m1_11639_23922# vss m1_12259_24224# vss nfet$150
Xpfet$145_2 vdd vdd m1_n5351_15778# m1_n4994_16080# pfet$145
Xpfet$150_0 vdd vdd vdd m1_33050_22344# m1_31535_22102# m1_31535_22102# pfet$150
Xnfet$178_3 m1_n9336_24346# m1_n9336_24346# vss vss m1_n9854_24542# vss nfet$178
Xpfet$144_11 vdd vdd m1_18705_21786# m1_18073_21786# pfet$144
Xnfet$157_8 m1_n7513_20152# vss m1_26676_16080# vss nfet$157
Xnfet$176_0 m1_n3822_20130# m1_n3822_20130# m1_n4485_20152# m1_n4485_20152# m1_n3724_20470#
+ vss nfet$176
Xnfet$183_1 m1_n2543_20130# m1_n2543_20130# m1_n5227_20152# m1_n5227_20152# m1_n2445_20470#
+ vss nfet$183
Xpfet$168_1 vdd m1_n8283_19850# m1_n8283_19850# m1_n8047_19550# m1_n8283_20611# m1_n8283_20611#
+ pfet$168
Xnfet$155_5 m1_965_15478# vss m1_8137_20152# vss nfet$155
Xnfet$153_28 m1_1933_17343# vss m1_2092_17836# vss nfet$153
Xnfet$153_17 m1_649_17714# vss m1_n2250_17343# vss nfet$153
Xnfet$153_39 m1_n3064_17714# vss m1_n3534_17714# vss nfet$153
Xnfet$162_6 m1_4637_21786# m1_4637_21786# vss vss m1_3475_21586# vss nfet$162
Xpfet$141_12 vdd m1_3989_15778# m1_3372_16080# m1_2092_17836# pfet$141
Xpfet$141_89 vdd vdd m1_22848_17343# m1_25747_17714# pfet$141
Xpfet$141_78 vdd vdd m1_13514_15478# sd4 pfet$141
Xpfet$141_67 vdd m1_22034_17714# vdd m1_23109_16202# pfet$141
Xpfet$141_23 vdd m1_5302_17714# vdd m1_6377_16202# pfet$141
Xpfet$141_34 vdd vdd m1_5761_16080# m1_n7513_20152# pfet$141
Xpfet$141_45 vdd vdd m1_9944_16080# m1_n7513_20152# pfet$141
Xpfet$141_56 vdd m1_n1278_18030# vdd m1_n2605_16080# pfet$141
Xnfet$153_2 m1_6275_17836# m1_7555_16080# m1_7088_18030# vss nfet$153
Xpfet$152_4 vdd m1_33174_24224# m1_34278_25658# m1_32193_25858# pfet$152
Xpfet$145_3 vdd vdd m1_n6657_17518# m1_n7247_17714# pfet$145
Xpfet$140_104 vdd m1_25912_25658# m1_26705_24542# m1_23964_25662# pfet$140
Xnfet$150_29 m1_15943_25858# vss m1_14556_21786# vss nfet$150
Xnfet$150_18 m1_7095_25858# vss m1_7232_25662# vss nfet$150
Xpfet$143_0 vdd m1_2590_19404# m1_2590_19404# m1_3458_19550# m1_n3534_17714# m1_n3534_17714#
+ pfet$143
Xnfet$178_4 m1_n4978_24224# m1_n4978_24224# m1_n10452_25858# m1_n10452_25858# m1_n4880_24542#
+ vss nfet$178
Xpfet$144_12 vdd vdd m1_16452_21590# m1_16322_21786# pfet$144
Xnfet$157_9 m1_n10452_25858# vss m1_27031_17343# vss nfet$157
Xnfet$169_0 m1_7198_15778# m1_7198_15778# m1_7088_18030# m1_7088_18030# m1_7324_17358#
+ vss nfet$169
Xnfet$176_1 m1_n1927_20274# m1_n1927_20274# vss vss m1_n2445_20470# vss nfet$176
Xpfet$168_2 vdd m1_n8283_20611# m1_n8283_20611# m1_n8047_22344# m1_n8145_21908# m1_n8145_21908#
+ pfet$168
Xnfet$153_29 m1_3372_16080# vss m1_3015_15778# vss nfet$153
Xnfet$153_18 m1_1119_17714# vss m1_649_17714# vss nfet$153
Xnfet$162_7 m1_488_21786# m1_488_21786# vss vss m1_n674_21586# vss nfet$162
Xnfet$155_6 m1_9015_17714# vss m1_12935_19550# vss nfet$155
Xpfet$141_79 vdd m1_15564_15778# m1_14743_16202# m1_14482_17343# pfet$141
Xpfet$141_68 vdd vdd m1_22034_17714# m1_22493_16080# pfet$141
Xpfet$141_13 vdd vdd m1_5148_15478# sd6 pfet$141
Xpfet$141_24 vdd m1_6377_16202# m1_5892_17518# m1_6275_17836# pfet$141
Xpfet$141_35 vdd vdd m1_9015_17714# m1_9485_17714# pfet$141
Xpfet$141_46 vdd vdd m1_n2250_17343# m1_649_17714# pfet$141
Xpfet$141_57 vdd m1_n1989_16202# m1_n2474_17518# m1_n2091_17836# pfet$141
Xpfet$166_10 vdd vdd m1_n10933_25858# fin pfet$166
Xnfet$153_3 m1_n7513_20152# vss m1_9944_16080# vss nfet$153
Xpfet$152_5 vdd m1_32817_25662# m1_32554_23922# m1_32330_25662# pfet$152
Xpfet$145_4 vdd vdd m1_n6433_17343# m1_n3534_17714# pfet$145
Xpfet$140_105 vdd vdd m1_30888_24542# m1_28492_25858# pfet$140
Xnfet$150_19 m1_7456_23922# vss m1_8076_24224# vss nfet$150
Xnfet$151_0 m1_n1133_21590# m1_n1133_21590# m1_354_22513# m1_354_22513# m1_n674_21586#
+ vss nfet$151
Xpfet$143_1 vdd vdd vdd m1_2822_19850# m1_4620_20152# m1_4620_20152# pfet$143
Xnfet$178_5 m1_n4362_24346# m1_n4362_24346# vss vss m1_n4880_24542# vss nfet$178
Xpfet$144_13 vdd vdd m1_15188_21786# m1_14556_21786# pfet$144
Xnfet$169_1 m1_5761_16080# m1_5761_16080# vss vss m1_7324_17358# vss nfet$169
Xnfet$176_2 m1_n3206_20274# m1_n3206_20274# vss vss m1_n3724_20470# vss nfet$176
Xnfet$153_19 m1_n7513_20152# vss m1_1578_16080# vss nfet$153
Xpfet$168_3 vdd vdd vdd m1_n8047_22344# m1_n8283_19850# m1_n8283_19850# pfet$168
Xnfet$162_8 m1_25739_21786# m1_25739_21786# vss vss m1_24577_21586# vss nfet$162
Xnfet$155_7 m1_5148_15478# vss m1_11654_20152# vss nfet$155
Xnfet$181_0 m1_n8283_20611# vss m1_n8283_19850# vss nfet$181
Xpfet$141_69 vdd vdd m1_20721_15778# m1_17851_17714# pfet$141
Xpfet$141_14 vdd vdd m1_2092_17836# m1_1933_17343# pfet$141
Xpfet$141_25 vdd vdd m1_1709_17518# m1_1119_17714# pfet$141
Xpfet$141_36 vdd vdd m1_6116_17343# m1_9015_17714# pfet$141
Xpfet$141_47 vdd m1_11738_16080# m1_11271_18030# m1_10299_17343# pfet$141
Xpfet$141_58 vdd vdd m1_n3534_17714# m1_n3064_17714# pfet$141
Xpfet$166_0 vdd vdd m1_n10796_25662# m1_n10933_25858# pfet$166
Xpfet$166_11 vdd vdd m1_n9336_24346# vss pfet$166
Xnfet$153_4 m1_10299_17343# m1_10560_16202# m1_10075_17518# vss nfet$153
Xpfet$152_6 vdd m1_34278_25658# m1_35071_24542# m1_32330_25662# pfet$152
Xpfet$145_5 vdd vdd m1_n6788_16080# m1_n7513_20152# pfet$145
Xpfet$140_106 vdd vdd m1_25107_21786# m1_28492_25858# pfet$140
Xnfet$151_1 m1_n1263_21786# m1_n1263_21786# m1_354_22513# m1_354_22513# m1_n42_21586#
+ vss nfet$151
Xpfet$143_2 vdd m1_2590_19404# m1_2590_19404# m1_2822_19850# m1_2384_19550# m1_2384_19550#
+ pfet$143
Xnfet$178_6 m1_n4978_24224# m1_n4978_24224# vss vss m1_n3415_25502# vss nfet$178
Xpfet$144_14 vdd vdd m1_19969_21590# m1_19839_21786# pfet$144
Xnfet$169_2 m1_9944_16080# m1_9944_16080# vss vss m1_11507_17358# vss nfet$169
Xnfet$176_3 m1_n6973_21481# m1_n6973_21481# m1_n6839_20152# m1_n6839_20152# m1_n6282_20470#
+ vss nfet$176
Xnfet$162_9 m1_25107_21786# m1_25107_21786# vss vss m1_23945_21586# vss nfet$162
Xnfet$155_8 m1_n7383_17599# vss m1_n1133_19550# vss nfet$155
Xpfet$141_15 vdd vdd m1_5302_17714# m1_5761_16080# pfet$141
Xpfet$141_26 vdd vdd m1_4832_17714# m1_5302_17714# pfet$141
Xpfet$141_37 vdd m1_7555_16080# m1_7088_18030# m1_6116_17343# pfet$141
Xpfet$141_48 vdd vdd m1_n3064_17714# m1_n2605_16080# pfet$141
Xnfet$181_1 m1_n7513_20152# m1_n8283_19850# vss vss nfet$181
Xpfet$141_59 vdd vdd m1_n2605_16080# m1_n7513_20152# pfet$141
Xpfet$166_1 vdd vdd m1_n10309_25662# m1_n10452_25858# pfet$166
Xnfet$174_0 m1_n10452_25858# m1_n10452_25858# m1_n7186_25858# m1_n7186_25858# m1_n6629_25502#
+ vss nfet$174
Xpfet$159_0 vdd m1_n4377_15778# m1_n4994_16080# m1_n6274_17836# pfet$159
Xpfet$166_12 vdd vdd m1_n7082_23622# m1_n8625_26174# pfet$166
Xpfet$152_7 vdd m1_32554_23922# m1_32818_24542# m1_32193_25858# pfet$152
Xnfet$153_5 m1_10458_17836# m1_11738_16080# m1_11271_18030# vss nfet$153
Xpfet$145_6 vdd vdd m1_n7383_17599# m1_n7247_17714# pfet$145
Xpfet$140_107 vdd m1_24309_25858# vdd m1_25912_25658# pfet$140
Xnfet$151_2 m1_9288_21786# m1_9288_21786# m1_9645_21447# m1_9645_21447# m1_10509_21586#
+ vss nfet$151
Xpfet$143_3 vdd vdd vdd m1_3458_19550# m1_n3218_15478# m1_n3218_15478# pfet$143
Xpfet$141_0 vdd vdd m1_12355_15778# m1_9485_17714# pfet$141
Xnfet$178_7 m1_n3541_23922# m1_n3541_23922# m1_n3651_26174# m1_n3651_26174# m1_n3415_25502#
+ vss nfet$178
Xpfet$144_15 vdd vdd m1_27003_21590# m1_26873_21786# pfet$144
Xnfet$169_3 m1_11381_15778# m1_11381_15778# m1_11271_18030# m1_11271_18030# m1_11507_17358#
+ vss nfet$169
Xnfet$176_4 m1_2590_19404# m1_2590_19404# vss vss m1_n2445_21430# vss nfet$176
Xnfet$155_9 m1_25747_17714# vss m1_27003_19550# vss nfet$155
Xnfet$167_0 m1_34093_22102# vss fout vss nfet$167
Xpfet$141_16 vdd vdd m1_3989_15778# m1_1119_17714# pfet$141
Xpfet$141_27 vdd m1_2194_16202# m1_1709_17518# m1_2092_17836# pfet$141
Xpfet$141_38 vdd vdd m1_7088_18030# m1_7198_15778# pfet$141
Xpfet$141_49 vdd m1_n194_15778# m1_n811_16080# m1_n2091_17836# pfet$141
Xnfet$181_2 m1_n8145_21908# vss m1_n8283_20611# vss nfet$181
Xnfet$174_1 m1_n6111_25858# m1_n6111_25858# vss vss m1_n6629_25502# vss nfet$174
Xpfet$159_1 vdd m1_n5351_15778# m1_n6172_16202# m1_n6433_17343# pfet$159
Xpfet$166_2 vdd vdd m1_n9952_24224# m1_n10572_23922# pfet$166
Xpfet$166_13 vdd vdd m1_n8055_24542# m1_n8625_26174# pfet$166
Xnfet$153_6 m1_6116_17343# vss m1_6275_17836# vss nfet$153
Xpfet$140_108 vdd vdd m1_25424_24346# m1_n7513_20152# pfet$140
Xpfet$145_7 vdd vdd m1_27190_17836# m1_27031_17343# pfet$145
Xpfet$171_0 vdd vdd vdd m1_n5019_19550# m1_n4485_20152# m1_n4485_20152# pfet$171
Xnfet$149_20 m1_21241_24346# m1_21241_24346# m1_20126_25858# m1_20126_25858# m1_22188_25502#
+ vss nfet$149
Xpfet$143_4 vdd m1_6107_19404# m1_6107_19404# m1_6339_19850# m1_5901_19550# m1_5901_19550#
+ pfet$143
Xnfet$151_3 m1_9418_21590# m1_9418_21590# m1_9645_21447# m1_9645_21447# m1_9877_21586#
+ vss nfet$151
Xnfet$151_10 m1_19839_21786# m1_19839_21786# m1_21456_22513# m1_21456_22513# m1_21060_21586#
+ vss nfet$151
Xpfet$141_1 vdd vdd m1_11381_15778# m1_11738_16080# pfet$141
Xpfet$144_16 vdd vdd m1_29256_21786# m1_28624_21786# pfet$144
Xnfet$176_5 m1_6107_19404# m1_6107_19404# m1_n5227_21418# m1_n5227_21418# m1_n2445_21430#
+ vss nfet$176
Xnfet$169_4 m1_10560_16202# m1_10560_16202# vss vss m1_10042_16398# vss nfet$169
Xpfet$141_17 vdd vdd m1_n2091_17836# m1_n2250_17343# pfet$141
Xnfet$181_3 m1_n8283_19850# m1_n8283_20611# vss vss nfet$181
Xpfet$141_28 vdd m1_2905_18030# vdd m1_1578_16080# pfet$141
Xpfet$141_39 vdd m1_7088_18030# vdd m1_5761_16080# pfet$141
Xpfet$159_2 vdd m1_n4994_16080# m1_n5461_18030# m1_n6433_17343# pfet$159
Xpfet$166_3 vdd vdd m1_n4978_24224# vss pfet$166
Xnfet$154_10 m1_21590_21786# vss m1_22222_21786# vss nfet$154
Xnfet$153_7 m1_9485_17714# vss m1_10075_17518# vss nfet$153
Xpfet$145_8 vdd vdd m1_28113_15778# m1_28470_16080# pfet$145
Xpfet$140_109 vdd m1_12259_24224# m1_13363_25658# m1_11278_25858# pfet$140
Xpfet$164_0 vdd vdd m1_n8625_26174# m1_n9336_24346# pfet$164
Xnfet$149_21 m1_28991_24224# m1_28991_24224# m1_28635_24542# m1_28635_24542# m1_29089_24542#
+ vss nfet$149
Xnfet$149_10 m1_17546_25658# m1_17546_25658# vss vss m1_18005_25502# vss nfet$149
Xpfet$143_5 vdd vdd vdd m1_n695_19850# m1_1103_20152# m1_1103_20152# pfet$143
Xnfet$151_4 m1_5901_21590# m1_5901_21590# m1_7388_22513# m1_7388_22513# m1_6360_21586#
+ vss nfet$151
Xnfet$151_11 m1_19969_21590# m1_19969_21590# m1_21456_22513# m1_21456_22513# m1_20428_21586#
+ vss nfet$151
Xpfet$141_2 vdd m1_12355_15778# m1_11738_16080# m1_10458_17836# pfet$141
Xpfet$144_17 vdd vdd m1_25739_21786# m1_25107_21786# pfet$144
Xnfet$162_10 m1_21590_21786# m1_21590_21786# vss vss m1_20428_21586# vss nfet$162
Xnfet$157_10 m1_26217_17714# vss m1_29087_15778# vss nfet$157
Xnfet$169_5 m1_9944_16080# m1_9944_16080# m1_9485_17714# m1_9485_17714# m1_10042_16398#
+ vss nfet$169
Xnfet$176_6 m1_n5764_21786# m1_n5764_21786# vss vss m1_n6282_21430# vss nfet$176
Xpfet$141_18 vdd m1_1119_17714# vdd m1_2194_16202# pfet$141
Xpfet$141_29 vdd vdd m1_1578_16080# m1_n7513_20152# pfet$141
Xpfet$159_3 vdd m1_n6172_16202# m1_n6657_17518# m1_n6274_17836# pfet$159
Xpfet$166_4 vdd vdd m1_n5571_25662# m1_n10452_25858# pfet$166
Xnfet$153_8 m1_7555_16080# vss m1_7198_15778# vss nfet$153
Xnfet$154_11 m1_18073_21786# vss m1_18705_21786# vss nfet$154
Xnfet$170_10 m1_9331_15478# m1_9331_15478# m1_n3822_21786# m1_n3822_21786# m1_13373_20470#
+ vss nfet$170
Xpfet$145_9 vdd vdd m1_29087_15778# m1_26217_17714# pfet$145
Xnfet$172_0 m1_n6274_17836# m1_n4994_16080# m1_n5461_18030# vss nfet$172
Xpfet$157_0 vdd m1_32818_20470# m1_32818_20470# m1_33050_19550# m1_30256_19792# m1_30256_19792#
+ pfet$157
Xpfet$164_1 vdd m1_n8625_26174# vdd m1_n8848_25658# pfet$164
Xnfet$149_22 m1_29607_24346# m1_29607_24346# vss vss m1_29089_24542# vss nfet$149
Xnfet$149_11 m1_16442_24224# m1_16442_24224# m1_16086_24542# m1_16086_24542# m1_16540_24542#
+ vss nfet$149
Xnfet$151_5 m1_2254_21786# m1_2254_21786# m1_3871_22513# m1_3871_22513# m1_3475_21586#
+ vss nfet$151
Xpfet$143_6 vdd vdd vdd m1_6339_19850# m1_8137_20152# m1_8137_20152# pfet$143
Xnfet$151_12 m1_16322_21786# m1_16322_21786# m1_17939_22513# m1_17939_22513# m1_17543_21586#
+ vss nfet$151
Xpfet$141_3 vdd m1_11381_15778# m1_10560_16202# m1_10299_17343# pfet$141
Xnfet$162_11 m1_22222_21786# m1_22222_21786# vss vss m1_21060_21586# vss nfet$162
Xnfet$157_11 m1_27031_17343# vss m1_27190_17836# vss nfet$157
Xnfet$169_6 m1_1578_16080# m1_1578_16080# vss vss m1_3141_17358# vss nfet$169
Xnfet$176_7 m1_n3822_21786# m1_n3822_21786# m1_n4485_21904# m1_n4485_21904# m1_n3724_21430#
+ vss nfet$176
Xpfet$159_4 vdd m1_28113_15778# m1_27292_16202# m1_27031_17343# pfet$159
Xpfet$141_19 vdd m1_3015_15778# m1_2194_16202# m1_1933_17343# pfet$141
Xpfet$166_5 vdd vdd m1_n4847_25662# m1_n10452_25858# pfet$166
Xnfet$153_9 sd5 vss m1_9331_15478# vss nfet$153
Xnfet$165_0 m1_31535_22102# m1_32818_21586# vss vss nfet$165
Xnfet$154_12 m1_14556_21786# vss m1_15188_21786# vss nfet$154
Xnfet$170_11 m1_15171_20152# m1_15171_20152# m1_n3822_21786# m1_n3822_21786# m1_14005_20470#
+ vss nfet$170
Xnfet$172_1 m1_n6433_17343# m1_n4377_15778# m1_n4994_16080# vss nfet$172
Xpfet$157_1 vdd vdd vdd m1_33050_19550# m1_31535_19792# m1_31535_19792# pfet$157
Xpfet$164_2 vdd m1_n3651_26174# vdd m1_n4978_24224# pfet$164
Xnfet$149_23 m1_25424_24346# m1_25424_24346# m1_24309_25858# m1_24309_25858# m1_26371_25502#
+ vss nfet$149
Xnfet$149_12 m1_17058_24346# m1_17058_24346# m1_15943_25858# m1_15943_25858# m1_18005_25502#
+ vss nfet$149
Xnfet$151_6 m1_2384_21590# m1_2384_21590# m1_3871_22513# m1_3871_22513# m1_2843_21586#
+ vss nfet$151
Xpfet$143_7 vdd vdd vdd m1_6975_19550# m1_965_15478# m1_965_15478# pfet$143
Xnfet$151_13 m1_16452_21590# m1_16452_21590# m1_17939_22513# m1_17939_22513# m1_16911_21586#
+ vss nfet$151
Xpfet$141_4 vdd m1_9485_17714# vdd m1_10560_16202# pfet$141
Xnfet$162_12 m1_18073_21786# m1_18073_21786# vss vss m1_16911_21586# vss nfet$162
Xnfet$157_12 m1_28470_16080# vss m1_28113_15778# vss nfet$157
Xnfet$169_7 m1_5761_16080# m1_5761_16080# m1_5302_17714# m1_5302_17714# m1_5859_16398#
+ vss nfet$169
Xnfet$176_8 m1_9624_19404# m1_9624_19404# vss vss m1_n3724_21430# vss nfet$176
Xpfet$166_6 vdd vdd m1_n4623_25487# fin pfet$166
Xpfet$159_5 vdd m1_29087_15778# m1_28470_16080# m1_27190_17836# pfet$159
Xnfet$154_13 m1_16322_21786# vss m1_16452_21590# vss nfet$154
Xnfet$170_12 m1_18688_20152# m1_18688_20152# m1_n1927_20274# m1_n1927_20274# m1_17522_20470#
+ vss nfet$170
Xnfet$172_2 m1_n6274_17836# m1_n5351_15778# m1_n6172_16202# vss nfet$172
Xpfet$157_2 vdd m1_32818_21586# m1_32818_21586# m1_33050_22344# m1_30256_22102# m1_30256_22102#
+ pfet$157
Xnfet$158_0 m1_n10452_25858# vss m1_n1271_25858# vss nfet$158
Xpfet$164_3 vdd vdd m1_n3651_26174# m1_n3541_23922# pfet$164
Xnfet$149_24 m1_30095_25658# m1_30095_25658# vss vss m1_30554_25502# vss nfet$149
Xnfet$149_13 m1_13363_25658# m1_13363_25658# vss vss m1_13822_25502# vss nfet$149
Xpfet$142_30 vdd vdd vdd m1_17539_22402# m1_16322_21786# m1_16322_21786# pfet$142
Xnfet$151_7 m1_5771_21786# m1_5771_21786# m1_7388_22513# m1_7388_22513# m1_6992_21586#
+ vss nfet$151
Xpfet$143_8 vdd m1_9624_19404# m1_9624_19404# m1_10492_19550# m1_4832_17714# m1_4832_17714#
+ pfet$143
Xpfet$162_0 vdd m1_n10309_25662# m1_n10572_23922# m1_n10796_25662# pfet$162
Xnfet$151_14 m1_12805_21786# m1_12805_21786# m1_14422_22513# m1_14422_22513# m1_14026_21586#
+ vss nfet$151
Xpfet$141_5 vdd m1_7198_15778# m1_6377_16202# m1_6116_17343# pfet$141
Xnfet$162_13 m1_18705_21786# m1_18705_21786# vss vss m1_17543_21586# vss nfet$162
Xnfet$157_13 m1_26217_17714# vss m1_25747_17714# vss nfet$157
Xnfet$169_8 m1_3015_15778# m1_3015_15778# m1_2905_18030# m1_2905_18030# m1_3141_17358#
+ vss nfet$169
Xnfet$176_9 m1_n6380_21786# m1_n6380_21786# m1_n6839_21786# m1_n6839_21786# m1_n6282_21430#
+ vss nfet$176
Xpfet$159_6 vdd m1_28470_16080# m1_28003_18030# m1_27031_17343# pfet$159
Xpfet$166_7 vdd vdd m1_n3541_23922# m1_n3184_24224# pfet$166
Xnfet$154_14 m1_19839_21786# vss m1_19969_21590# vss nfet$154
Xnfet$170_13 m1_13514_15478# m1_13514_15478# m1_n1927_20274# m1_n1927_20274# m1_16890_20470#
+ vss nfet$170
Xnfet$172_3 m1_n6433_17343# m1_n6172_16202# m1_n6657_17518# vss nfet$172
Xnfet$158_1 m1_n789_25858# vss m1_n647_25662# vss nfet$158
Xpfet$164_4 vdd m1_n10452_25858# vdd m1_n4362_24346# pfet$164
Xpfet$142_31 vdd vdd vdd m1_27462_22102# m1_27003_21590# m1_27003_21590# pfet$142
Xnfet$149_14 m1_12875_24346# m1_12875_24346# m1_11760_25858# m1_11760_25858# m1_13822_25502#
+ vss nfet$149
Xpfet$142_20 vdd vdd vdd m1_20428_22102# m1_19969_21590# m1_19969_21590# pfet$142
Xnfet$149_25 m1_29607_24346# m1_29607_24346# m1_28492_25858# m1_28492_25858# m1_30554_25502#
+ vss nfet$149
Xnfet$151_8 m1_23486_21590# m1_23486_21590# m1_24973_22513# m1_24973_22513# m1_23945_21586#
+ vss nfet$151
Xnfet$170_0 m1_4620_20152# m1_4620_20152# m1_2590_19404# m1_2590_19404# m1_3454_20470#
+ vss nfet$170
Xpfet$143_9 vdd m1_9624_19404# m1_9624_19404# m1_9856_19850# m1_9418_19550# m1_9418_19550#
+ pfet$143
Xpfet$155_0 vdd vdd vdd m1_36073_22344# define define pfet$155
Xpfet$162_1 vdd m1_n9952_24224# m1_n8848_25658# m1_n10933_25858# pfet$162
Xnfet$151_15 m1_26873_21786# m1_26873_21786# m1_28490_22513# m1_28490_22513# m1_28094_21586#
+ vss nfet$151
Xpfet$141_6 vdd vdd m1_7198_15778# m1_7555_16080# pfet$141
Xnfet$162_14 m1_15188_21786# m1_15188_21786# vss vss m1_14026_21586# vss nfet$162
.ends

.subckt pfet$208 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$206 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$221 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt nfet$219 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$209 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$207 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$222 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$220 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt asc_drive_buffer vss in vdd out
Xpfet$208_0 vdd vdd m1_4002_n1060# m1_3466_n454# pfet$208
Xpfet$206_0 out out m1_4274_n1060# vdd m1_4274_n1060# out vdd vdd m1_4274_n1060# out
+ m1_4274_n1060# m1_4274_n1060# out m1_4274_n1060# vdd m1_4274_n1060# vdd m1_4274_n1060#
+ pfet$206
Xnfet$221_0 m1_3466_n454# vss m1_4002_n1060# vss nfet$221
Xnfet$219_0 m1_4274_n1060# vss m1_4002_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ m1_4274_n1060# vss m1_4002_n1060# vss nfet$219
Xpfet$209_0 vdd vdd m1_3466_n454# in pfet$209
Xpfet$207_0 m1_4274_n1060# vdd vdd m1_4274_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ vdd m1_4002_n1060# m1_4002_n1060# pfet$207
Xnfet$222_0 in vss m1_3466_n454# vss nfet$222
Xnfet$220_0 out out vss m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# m1_4274_n1060#
+ m1_4274_n1060# out m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# vss vss
+ nfet$220
.ends

.subckt nfet$213 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$199 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$212 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$200 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt xp_3_1_MUX$1 S0 S1 VDD VSS OUT_1 C_1 B_1 A_1
Xnfet$213_0 S1 VSS m1_n432_n1290# VSS nfet$213
Xnfet$213_1 S0 VSS m1_n432_458# VSS nfet$213
Xpfet$199_0 VDD A_1 m1_239_n318# m1_n432_458# pfet$199
Xpfet$199_1 VDD C_1 OUT_1 S1 pfet$199
Xpfet$199_2 VDD B_1 m1_239_n318# S0 pfet$199
Xpfet$199_3 VDD m1_239_n318# OUT_1 m1_n432_n1290# pfet$199
Xnfet$212_0 m1_n432_n1290# C_1 OUT_1 VSS nfet$212
Xnfet$212_1 m1_n432_458# B_1 m1_239_n318# VSS nfet$212
Xnfet$212_2 S1 m1_239_n318# OUT_1 VSS nfet$212
Xnfet$212_3 S0 A_1 m1_239_n318# VSS nfet$212
Xpfet$200_0 VDD VDD m1_n432_n1290# S1 pfet$200
Xpfet$200_1 VDD VDD m1_n432_458# S0 pfet$200
.ends

.subckt nfet$193 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$183 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$181 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$196 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$179 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$194 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$192 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$182 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$180 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$195 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt asc_hysteresis_buffer$2 vss in vdd out
Xnfet$193_0 m1_348_648# vss m1_884_42# vss nfet$193
Xpfet$183_0 vdd vdd m1_884_42# m1_1156_42# pfet$183
Xpfet$181_0 vdd vdd m1_348_648# in pfet$181
Xnfet$196_0 m1_1156_42# vss m1_884_42# vss nfet$196
Xpfet$179_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd
+ m1_884_42# m1_884_42# pfet$179
Xnfet$194_0 in vss m1_348_648# vss nfet$194
Xnfet$192_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$192
Xpfet$182_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$182
Xpfet$180_0 vdd vdd m1_884_42# m1_348_648# pfet$180
Xnfet$195_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$195
.ends

.subckt nfet$197 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$189 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$187 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$185 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$192 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$206 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$190 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$211 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$204 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$202 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$197 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$200 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt nfet$198 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$195 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=0.78p ps=3.52u w=3u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.78p pd=3.52u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$188 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$209 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$193 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt pfet$186 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$207 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$191 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt pfet$184 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$205 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$210 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$203 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$198 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$201 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt nfet$199 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$196 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$194 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$208 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_lock_detector_20250826 ref vdd div vss lock
Xnfet$197_5 m1_8596_7868# m1_8596_7868# vss m1_7448_4493# m1_7448_4493# m1_8596_7868#
+ vss m1_7448_4493# m1_7448_4493# m1_7448_4493# m1_8596_7868# m1_7448_4493# m1_7448_4493#
+ m1_8596_7868# vss m1_7448_4493# vss vss nfet$197
Xpfet$189_6 vdd m1_16599_5522# m1_17703_6956# m1_15618_7156# pfet$189
Xpfet$187_3 m1_n940_n340# vdd vdd m1_n940_n340# m1_n1212_n340# m1_n1212_n340# m1_n940_n340#
+ vdd m1_n1212_n340# m1_n1212_n340# pfet$187
Xpfet$185_0 vdd vdd m1_7176_n340# m1_6640_1478# pfet$185
Xpfet$192_1 m1_n7214_4493# vdd vdd m1_n7214_4493# m1_n7486_4493# m1_n7486_4493# m1_n7214_4493#
+ vdd m1_n7486_4493# m1_n7486_4493# pfet$192
Xnfet$197_6 m1_208_7868# m1_208_7868# vss m1_n940_4493# m1_n940_4493# m1_208_7868#
+ vss m1_n940_4493# m1_n940_4493# m1_n940_4493# m1_208_7868# m1_n940_4493# m1_n940_4493#
+ m1_208_7868# vss m1_n940_4493# vss vss nfet$197
Xpfet$189_7 vdd m1_16242_6960# m1_15979_5220# m1_15755_6960# pfet$189
Xpfet$187_4 m1_n940_4493# vdd vdd m1_n940_4493# m1_n1212_4493# m1_n1212_4493# m1_n940_4493#
+ vdd m1_n1212_4493# m1_n1212_4493# pfet$187
Xnfet$206_0 m1_15979_2344# vss m1_16599_2028# vss nfet$206
Xpfet$185_1 vdd vdd m1_11370_n340# m1_10834_1478# pfet$185
Xpfet$192_2 m1_n15602_4493# vdd vdd m1_n15602_4493# m1_n15874_4493# m1_n15874_4493#
+ m1_n15602_4493# vdd m1_n15874_4493# m1_n15874_4493# pfet$192
Xnfet$197_7 m1_4402_7868# m1_4402_7868# vss m1_3254_4493# m1_3254_4493# m1_4402_7868#
+ vss m1_3254_4493# m1_3254_4493# m1_3254_4493# m1_4402_7868# m1_3254_4493# m1_3254_4493#
+ m1_4402_7868# vss m1_3254_4493# vss vss nfet$197
Xpfet$187_5 m1_11642_4493# vdd vdd m1_11642_4493# m1_11370_4493# m1_11370_4493# m1_11642_4493#
+ vdd m1_11370_4493# m1_11370_4493# pfet$187
Xpfet$185_2 vdd vdd m1_2982_n340# m1_2446_1478# pfet$185
Xpfet$190_0 vdd m1_17926_34# vdd m1_17703_788# pfet$190
Xnfet$206_1 m1_15618_394# vss m1_15755_n208# vss nfet$206
Xpfet$187_6 m1_3254_4493# vdd vdd m1_3254_4493# m1_2982_4493# m1_2982_4493# m1_3254_4493#
+ vdd m1_2982_4493# m1_2982_4493# pfet$187
Xpfet$190_1 vdd vdd m1_17926_34# m1_17215_2028# pfet$190
Xnfet$206_2 m1_n2336_5099# vss m1_16242_n208# vss nfet$206
Xpfet$185_3 vdd vdd m1_n1212_n340# m1_n1748_1478# pfet$185
Xnfet$211_0 m1_19675_2344# vss lock vss nfet$211
Xpfet$187_7 m1_7448_4493# vdd vdd m1_7448_4493# m1_7176_4493# m1_7176_4493# m1_7448_4493#
+ vdd m1_7176_4493# m1_7176_4493# pfet$187
Xpfet$185_4 vdd vdd m1_n1212_4493# m1_n1748_5099# pfet$185
Xnfet$204_0 m1_15755_n208# m1_16599_2028# m1_17703_788# vss nfet$204
Xpfet$190_2 vdd m1_16243_1828# vdd m1_17215_2028# pfet$190
Xnfet$206_3 m1_17926_34# vss m1_18496_1828# vss nfet$206
Xpfet$185_5 vdd vdd m1_2982_4493# m1_2446_5099# pfet$185
Xpfet$190_3 vdd vdd m1_16243_1828# m1_16599_2028# pfet$190
Xnfet$206_4 m1_12790_n340# vss m1_15618_394# vss nfet$206
Xnfet$204_1 m1_15618_394# m1_16242_n208# m1_15979_2344# vss nfet$204
Xpfet$185_6 vdd vdd m1_7176_4493# m1_6640_5099# pfet$185
Xnfet$204_2 m1_15618_394# m1_17703_788# m1_18496_1828# vss nfet$204
Xnfet$206_5 vss vss m1_17215_2028# vss nfet$206
Xpfet$190_4 vdd m1_16243_5840# vdd m1_17215_5644# pfet$190
Xpfet$185_7 vdd vdd m1_11370_4493# m1_10834_5099# pfet$185
Xnfet$206_6 m1_17926_34# vss m1_19469_1832# vss nfet$206
Xpfet$190_5 vdd vdd m1_16243_5840# m1_16599_5522# pfet$190
Xnfet$204_3 m1_15755_n208# m1_15979_2344# m1_16243_1828# vss nfet$204
Xnfet$202_0 m1_n7214_4493# vss m1_n7486_4493# m1_n7486_4493# m1_n7486_4493# m1_n7214_4493#
+ m1_n7214_4493# vss m1_n7486_4493# vss nfet$202
Xpfet$190_6 vdd m1_17926_7472# vdd m1_17703_6956# pfet$190
Xnfet$206_7 vss vss m1_17215_5644# vss nfet$206
Xnfet$202_1 m1_n15602_4493# vss m1_n15874_4493# m1_n15874_4493# m1_n15874_4493# m1_n15602_4493#
+ m1_n15602_4493# vss m1_n15874_4493# vss nfet$202
Xnfet$204_4 m1_15618_7156# m1_17703_6956# m1_18496_5840# vss nfet$204
Xnfet$206_8 m1_17926_7472# vss m1_19469_4920# vss nfet$206
Xpfet$197_0 vdd m1_19675_2344# vdd m1_19469_1832# pfet$197
Xpfet$190_7 vdd vdd m1_17926_7472# m1_17215_5644# pfet$190
Xnfet$204_5 m1_15755_6960# m1_15979_5220# m1_16243_5840# vss nfet$204
Xnfet$202_2 m1_n11408_4493# vss m1_n11680_4493# m1_n11680_4493# m1_n11680_4493# m1_n11408_4493#
+ m1_n11408_4493# vss m1_n11680_4493# vss nfet$202
Xnfet$206_9 m1_17926_7472# vss m1_18496_5840# vss nfet$206
Xpfet$197_1 vdd vdd m1_19675_2344# m1_19469_4920# pfet$197
Xnfet$204_6 m1_15618_7156# m1_16242_6960# m1_15979_5220# vss nfet$204
Xnfet$200_0 m1_n6066_7868# m1_n6066_7868# vss m1_n7214_4493# m1_n7214_4493# m1_n6066_7868#
+ vss m1_n7214_4493# m1_n7214_4493# m1_n7214_4493# m1_n6066_7868# m1_n7214_4493# m1_n7214_4493#
+ m1_n6066_7868# vss m1_n7214_4493# vss vss nfet$200
Xnfet$198_0 m1_10834_1478# vss m1_11370_n340# vss nfet$198
Xnfet$204_7 m1_15755_6960# m1_16599_5522# m1_17703_6956# vss nfet$204
Xnfet$200_1 m1_n14454_7868# m1_n14454_7868# vss m1_n15602_4493# m1_n15602_4493# m1_n14454_7868#
+ vss m1_n15602_4493# m1_n15602_4493# m1_n15602_4493# m1_n14454_7868# m1_n15602_4493#
+ m1_n15602_4493# m1_n14454_7868# vss m1_n15602_4493# vss vss nfet$200
Xnfet$198_1 m1_2446_1478# vss m1_2982_n340# vss nfet$198
Xpfet$195_0 vdd vdd vdd m1_n3798_6028# div div pfet$195
Xnfet$200_2 m1_n10260_7868# m1_n10260_7868# vss m1_n11408_4493# m1_n11408_4493# m1_n10260_7868#
+ vss m1_n11408_4493# m1_n11408_4493# m1_n11408_4493# m1_n10260_7868# m1_n11408_4493#
+ m1_n11408_4493# m1_n10260_7868# vss m1_n11408_4493# vss vss nfet$200
Xnfet$198_2 m1_6640_1478# vss m1_7176_n340# vss nfet$198
Xpfet$188_0 vdd vdd m1_16599_2028# m1_15979_2344# pfet$188
Xpfet$195_1 vdd m1_n4030_5270# m1_n4030_5270# m1_n3798_6028# m1_n6066_7868# m1_n6066_7868#
+ pfet$195
Xnfet$198_3 m1_n1748_1478# vss m1_n1212_n340# vss nfet$198
Xpfet$188_1 vdd vdd m1_16242_n208# m1_n2336_5099# pfet$188
Xnfet$209_0 m1_n4030_5270# vss m1_n2336_5099# vss nfet$209
Xnfet$198_4 m1_10834_5099# vss m1_11370_4493# vss nfet$198
Xpfet$188_2 vdd vdd m1_15755_n208# m1_15618_394# pfet$188
Xpfet$193_0 vdd vdd m1_n11680_4493# m1_n12216_5099# pfet$193
Xnfet$198_5 m1_6640_5099# vss m1_7176_4493# vss nfet$198
Xpfet$188_3 vdd vdd m1_18496_1828# m1_17926_34# pfet$188
Xpfet$186_0 m1_8596_n340# m1_8596_n340# m1_7448_n340# vdd m1_7448_n340# m1_8596_n340#
+ vdd vdd m1_7448_n340# m1_8596_n340# m1_7448_n340# m1_7448_n340# m1_8596_n340# m1_7448_n340#
+ vdd m1_7448_n340# vdd m1_7448_n340# pfet$186
Xpfet$193_1 vdd vdd m1_n7486_4493# m1_n8022_5099# pfet$193
Xnfet$198_6 m1_n1748_5099# vss m1_n1212_4493# vss nfet$198
Xpfet$188_4 vdd vdd m1_15618_394# m1_12790_n340# pfet$188
Xpfet$186_1 m1_12790_n340# m1_12790_n340# m1_11642_n340# vdd m1_11642_n340# m1_12790_n340#
+ vdd vdd m1_11642_n340# m1_12790_n340# m1_11642_n340# m1_11642_n340# m1_12790_n340#
+ m1_11642_n340# vdd m1_11642_n340# vdd m1_11642_n340# pfet$186
Xnfet$207_0 m1_n14454_7868# vss m1_n12216_5099# vss nfet$207
Xpfet$193_2 vdd vdd m1_n15874_4493# m1_n16410_5099# pfet$193
Xnfet$198_7 m1_2446_5099# vss m1_2982_4493# vss nfet$198
Xpfet$188_5 vdd vdd m1_17215_2028# vss pfet$188
Xpfet$186_2 m1_4402_n340# m1_4402_n340# m1_3254_n340# vdd m1_3254_n340# m1_4402_n340#
+ vdd vdd m1_3254_n340# m1_4402_n340# m1_3254_n340# m1_3254_n340# m1_4402_n340# m1_3254_n340#
+ vdd m1_3254_n340# vdd m1_3254_n340# pfet$186
Xnfet$207_1 div vss m1_n16410_5099# vss nfet$207
Xpfet$191_0 m1_n10260_7868# m1_n10260_7868# m1_n11408_4493# vdd m1_n11408_4493# m1_n10260_7868#
+ vdd vdd m1_n11408_4493# m1_n10260_7868# m1_n11408_4493# m1_n11408_4493# m1_n10260_7868#
+ m1_n11408_4493# vdd m1_n11408_4493# vdd m1_n11408_4493# pfet$191
Xpfet$188_6 vdd vdd m1_19469_1832# m1_17926_34# pfet$188
Xpfet$186_3 m1_208_n340# m1_208_n340# m1_n940_n340# vdd m1_n940_n340# m1_208_n340#
+ vdd vdd m1_n940_n340# m1_208_n340# m1_n940_n340# m1_n940_n340# m1_208_n340# m1_n940_n340#
+ vdd m1_n940_n340# vdd m1_n940_n340# pfet$186
Xnfet$207_2 m1_n10260_7868# vss m1_n8022_5099# vss nfet$207
Xpfet$184_0 vdd vdd m1_6640_1478# m1_4402_n340# pfet$184
Xpfet$191_1 m1_n6066_7868# m1_n6066_7868# m1_n7214_4493# vdd m1_n7214_4493# m1_n6066_7868#
+ vdd vdd m1_n7214_4493# m1_n6066_7868# m1_n7214_4493# m1_n7214_4493# m1_n6066_7868#
+ m1_n7214_4493# vdd m1_n7214_4493# vdd m1_n7214_4493# pfet$191
Xpfet$188_7 vdd vdd m1_17215_5644# vss pfet$188
Xpfet$184_1 vdd vdd m1_10834_1478# m1_8596_n340# pfet$184
Xpfet$186_4 m1_208_7868# m1_208_7868# m1_n940_4493# vdd m1_n940_4493# m1_208_7868#
+ vdd vdd m1_n940_4493# m1_208_7868# m1_n940_4493# m1_n940_4493# m1_208_7868# m1_n940_4493#
+ vdd m1_n940_4493# vdd m1_n940_4493# pfet$186
Xpfet$191_2 m1_n14454_7868# m1_n14454_7868# m1_n15602_4493# vdd m1_n15602_4493# m1_n14454_7868#
+ vdd vdd m1_n15602_4493# m1_n14454_7868# m1_n15602_4493# m1_n15602_4493# m1_n14454_7868#
+ m1_n15602_4493# vdd m1_n15602_4493# vdd m1_n15602_4493# pfet$191
Xnfet$205_0 m1_17215_2028# m1_17215_2028# m1_17926_34# m1_17926_34# m1_18162_712#
+ vss nfet$205
Xpfet$188_8 vdd vdd m1_19469_4920# m1_17926_7472# pfet$188
Xpfet$186_5 m1_12790_7868# m1_12790_7868# m1_11642_4493# vdd m1_11642_4493# m1_12790_7868#
+ vdd vdd m1_11642_4493# m1_12790_7868# m1_11642_4493# m1_11642_4493# m1_12790_7868#
+ m1_11642_4493# vdd m1_11642_4493# vdd m1_11642_4493# pfet$186
Xnfet$205_1 m1_17703_788# m1_17703_788# vss vss m1_18162_712# vss nfet$205
Xpfet$184_2 vdd vdd m1_n1748_1478# ref pfet$184
Xpfet$188_9 vdd vdd m1_18496_5840# m1_17926_7472# pfet$188
Xpfet$186_6 m1_4402_7868# m1_4402_7868# m1_3254_4493# vdd m1_3254_4493# m1_4402_7868#
+ vdd vdd m1_3254_4493# m1_4402_7868# m1_3254_4493# m1_3254_4493# m1_4402_7868# m1_3254_4493#
+ vdd m1_3254_4493# vdd m1_3254_4493# pfet$186
Xpfet$184_3 vdd vdd m1_n1748_5099# m1_n2336_5099# pfet$184
Xnfet$205_2 m1_16599_2028# m1_16599_2028# m1_16243_1828# m1_16243_1828# m1_16697_1672#
+ vss nfet$205
Xnfet$210_0 m1_19469_4920# m1_19469_4920# m1_19675_2344# m1_19675_2344# m1_19911_1672#
+ vss nfet$210
Xpfet$186_7 m1_8596_7868# m1_8596_7868# m1_7448_4493# vdd m1_7448_4493# m1_8596_7868#
+ vdd vdd m1_7448_4493# m1_8596_7868# m1_7448_4493# m1_7448_4493# m1_8596_7868# m1_7448_4493#
+ vdd m1_7448_4493# vdd m1_7448_4493# pfet$186
Xpfet$184_4 vdd vdd m1_6640_5099# m1_4402_7868# pfet$184
Xnfet$205_3 m1_17215_2028# m1_17215_2028# vss vss m1_16697_1672# vss nfet$205
Xnfet$203_0 m1_8596_n340# vss m1_10834_1478# vss nfet$203
Xnfet$210_1 m1_19469_1832# m1_19469_1832# vss vss m1_19911_1672# vss nfet$210
Xpfet$184_5 vdd vdd m1_10834_5099# m1_8596_7868# pfet$184
Xnfet$205_4 m1_17215_5644# m1_17215_5644# vss vss m1_16697_5840# vss nfet$205
Xnfet$203_1 m1_4402_n340# vss m1_6640_1478# vss nfet$203
Xpfet$184_6 vdd vdd m1_2446_5099# m1_208_7868# pfet$184
Xnfet$205_5 m1_16599_5522# m1_16599_5522# m1_16243_5840# m1_16243_5840# m1_16697_5840#
+ vss nfet$205
Xpfet$198_0 vdd vdd lock m1_19675_2344# pfet$198
Xnfet$203_2 ref vss m1_n1748_1478# vss nfet$203
Xpfet$184_7 vdd vdd m1_2446_1478# m1_208_n340# pfet$184
Xnfet$205_6 m1_17215_5644# m1_17215_5644# m1_17926_7472# m1_17926_7472# m1_18162_6800#
+ vss nfet$205
Xnfet$201_0 m1_n8022_5099# vss m1_n7486_4493# vss nfet$201
Xnfet$203_3 m1_n2336_5099# vss m1_n1748_5099# vss nfet$203
Xnfet$199_0 m1_3254_n340# vss m1_2982_n340# m1_2982_n340# m1_2982_n340# m1_3254_n340#
+ m1_3254_n340# vss m1_2982_n340# vss nfet$199
Xnfet$205_7 m1_17703_6956# m1_17703_6956# vss vss m1_18162_6800# vss nfet$205
Xnfet$206_10 m1_12790_7868# vss m1_15618_7156# vss nfet$206
Xnfet$203_4 m1_8596_7868# vss m1_10834_5099# vss nfet$203
Xnfet$201_1 m1_n16410_5099# vss m1_n15874_4493# vss nfet$201
Xnfet$199_1 m1_7448_n340# vss m1_7176_n340# m1_7176_n340# m1_7176_n340# m1_7448_n340#
+ m1_7448_n340# vss m1_7176_n340# vss nfet$199
Xnfet$206_11 m1_15979_5220# vss m1_16599_5522# vss nfet$206
Xpfet$196_0 vdd vdd m1_n2336_5099# m1_n4030_5270# pfet$196
Xnfet$201_2 m1_n12216_5099# vss m1_n11680_4493# vss nfet$201
Xnfet$203_5 m1_4402_7868# vss m1_6640_5099# vss nfet$203
Xpfet$188_10 vdd vdd m1_15618_7156# m1_12790_7868# pfet$188
Xnfet$206_12 m1_15618_7156# vss m1_15755_6960# vss nfet$206
Xpfet$189_0 vdd m1_16599_2028# m1_17703_788# m1_15618_394# pfet$189
Xnfet$199_2 m1_11642_n340# vss m1_11370_n340# m1_11370_n340# m1_11370_n340# m1_11642_n340#
+ m1_11642_n340# vss m1_11370_n340# vss nfet$199
Xnfet$203_6 m1_208_n340# vss m1_2446_1478# vss nfet$203
Xpfet$188_11 vdd vdd m1_16599_5522# m1_15979_5220# pfet$188
Xnfet$199_3 m1_n940_n340# vss m1_n1212_n340# m1_n1212_n340# m1_n1212_n340# m1_n940_n340#
+ m1_n940_n340# vss m1_n1212_n340# vss nfet$199
Xnfet$206_13 ref vss m1_16242_6960# vss nfet$206
Xpfet$189_1 vdd m1_16242_n208# m1_15979_2344# m1_15755_n208# pfet$189
Xnfet$197_0 m1_8596_n340# m1_8596_n340# vss m1_7448_n340# m1_7448_n340# m1_8596_n340#
+ vss m1_7448_n340# m1_7448_n340# m1_7448_n340# m1_8596_n340# m1_7448_n340# m1_7448_n340#
+ m1_8596_n340# vss m1_7448_n340# vss vss nfet$197
Xnfet$203_7 m1_208_7868# vss m1_2446_5099# vss nfet$203
Xpfet$188_12 vdd vdd m1_16242_6960# ref pfet$188
Xnfet$199_4 m1_11642_4493# vss m1_11370_4493# m1_11370_4493# m1_11370_4493# m1_11642_4493#
+ m1_11642_4493# vss m1_11370_4493# vss nfet$199
Xnfet$197_1 m1_4402_n340# m1_4402_n340# vss m1_3254_n340# m1_3254_n340# m1_4402_n340#
+ vss m1_3254_n340# m1_3254_n340# m1_3254_n340# m1_4402_n340# m1_3254_n340# m1_3254_n340#
+ m1_4402_n340# vss m1_3254_n340# vss vss nfet$197
Xpfet$189_2 vdd m1_15979_2344# m1_16243_1828# m1_15618_394# pfet$189
Xpfet$194_0 vdd vdd m1_n8022_5099# m1_n10260_7868# pfet$194
Xnfet$199_5 m1_7448_4493# vss m1_7176_4493# m1_7176_4493# m1_7176_4493# m1_7448_4493#
+ m1_7448_4493# vss m1_7176_4493# vss nfet$199
Xpfet$188_13 vdd vdd m1_15755_6960# m1_15618_7156# pfet$188
Xnfet$197_2 m1_12790_n340# m1_12790_n340# vss m1_11642_n340# m1_11642_n340# m1_12790_n340#
+ vss m1_11642_n340# m1_11642_n340# m1_11642_n340# m1_12790_n340# m1_11642_n340# m1_11642_n340#
+ m1_12790_n340# vss m1_11642_n340# vss vss nfet$197
Xpfet$189_3 vdd m1_17703_788# m1_18496_1828# m1_15755_n208# pfet$189
Xpfet$187_0 m1_7448_n340# vdd vdd m1_7448_n340# m1_7176_n340# m1_7176_n340# m1_7448_n340#
+ vdd m1_7176_n340# m1_7176_n340# pfet$187
Xpfet$194_1 vdd vdd m1_n16410_5099# div pfet$194
Xnfet$199_6 m1_n940_4493# vss m1_n1212_4493# m1_n1212_4493# m1_n1212_4493# m1_n940_4493#
+ m1_n940_4493# vss m1_n1212_4493# vss nfet$199
Xnfet$197_3 m1_208_n340# m1_208_n340# vss m1_n940_n340# m1_n940_n340# m1_208_n340#
+ vss m1_n940_n340# m1_n940_n340# m1_n940_n340# m1_208_n340# m1_n940_n340# m1_n940_n340#
+ m1_208_n340# vss m1_n940_n340# vss vss nfet$197
Xpfet$189_4 vdd m1_17703_6956# m1_18496_5840# m1_15755_6960# pfet$189
Xpfet$187_1 m1_11642_n340# vdd vdd m1_11642_n340# m1_11370_n340# m1_11370_n340# m1_11642_n340#
+ vdd m1_11370_n340# m1_11370_n340# pfet$187
Xpfet$194_2 vdd vdd m1_n12216_5099# m1_n14454_7868# pfet$194
Xnfet$208_0 div m1_n4030_5270# vss vss nfet$208
Xnfet$199_7 m1_3254_4493# vss m1_2982_4493# m1_2982_4493# m1_2982_4493# m1_3254_4493#
+ m1_3254_4493# vss m1_2982_4493# vss nfet$199
Xnfet$197_4 m1_12790_7868# m1_12790_7868# vss m1_11642_4493# m1_11642_4493# m1_12790_7868#
+ vss m1_11642_4493# m1_11642_4493# m1_11642_4493# m1_12790_7868# m1_11642_4493# m1_11642_4493#
+ m1_12790_7868# vss m1_11642_4493# vss vss nfet$197
Xpfet$189_5 vdd m1_15979_5220# m1_16243_5840# m1_15618_7156# pfet$189
Xpfet$187_2 m1_3254_n340# vdd vdd m1_3254_n340# m1_2982_n340# m1_2982_n340# m1_3254_n340#
+ vdd m1_2982_n340# m1_2982_n340# pfet$187
Xnfet$208_1 m1_n6066_7868# vss m1_n4030_5270# vss nfet$208
Xpfet$192_0 m1_n11408_4493# vdd vdd m1_n11408_4493# m1_n11680_4493# m1_n11680_4493#
+ m1_n11408_4493# vdd m1_n11680_4493# m1_n11680_4493# pfet$192
.ends

.subckt asc_dual_psd_def_20250809$1 vdd vss pd1 pd2 pd3 pd4 pd5 pd6 pd7 pd8 pd9 fout
+ sd1 sd2 sd3 sd4 sd5 sd6 sd7 sd8 sd9 fin define
Xnfet$169_9 m1_2194_16202# m1_2194_16202# vss vss m1_1676_16398# vss nfet$169
Xpfet$159_7 vdd m1_27292_16202# m1_26807_17518# m1_27190_17836# pfet$159
Xpfet$166_8 vdd vdd m1_n2567_23922# m1_n7320_25516# pfet$166
Xnfet$154_15 m1_28624_21786# vss m1_29256_21786# vss nfet$154
Xnfet$170_14 m1_22205_20152# m1_22205_20152# m1_n2543_20130# m1_n2543_20130# m1_21039_20470#
+ vss nfet$170
Xnfet$172_4 m1_27031_17343# m1_27292_16202# m1_26807_17518# vss nfet$172
Xnfet$158_2 m1_n1271_25858# vss m1_n1134_25662# vss nfet$158
Xpfet$142_32 vdd m1_28490_22513# m1_28490_22513# m1_28090_22402# m1_28624_21786# m1_28624_21786#
+ pfet$142
Xpfet$142_21 vdd vdd vdd m1_21056_22402# m1_19839_21786# m1_19839_21786# pfet$142
Xpfet$164_5 vdd vdd m1_n10308_24542# m1_n9952_24224# pfet$164
Xpfet$142_10 vdd m1_3871_22513# m1_3871_22513# m1_2843_22102# m1_4637_21786# m1_4637_21786#
+ pfet$142
Xnfet$149_26 m1_25912_25658# m1_25912_25658# vss vss m1_26371_25502# vss nfet$149
Xnfet$149_15 m1_25424_24346# m1_25424_24346# vss vss m1_24906_24542# vss nfet$149
Xnfet$151_9 m1_23356_21786# m1_23356_21786# m1_24973_22513# m1_24973_22513# m1_24577_21586#
+ vss nfet$151
Xnfet$170_1 m1_1103_20152# m1_1103_20152# m1_n927_19404# m1_n927_19404# m1_n63_20470#
+ vss nfet$170
Xpfet$155_1 vdd m1_35837_22102# m1_35837_22102# m1_36073_22344# fout fout pfet$155
Xnfet$163_0 m1_21456_22513# m1_21456_22513# m1_30256_19792# m1_30256_19792# m1_30492_20470#
+ vss nfet$163
Xpfet$162_2 vdd m1_n4362_24346# m1_n4847_25662# m1_n4464_25980# pfet$162
Xpfet$148_0 vdd vdd m1_n647_25662# m1_n789_25858# pfet$148
Xnfet$151_16 m1_27003_21590# m1_27003_21590# m1_28490_22513# m1_28490_22513# m1_27462_21586#
+ vss nfet$151
Xpfet$141_7 vdd vdd m1_6275_17836# m1_6116_17343# pfet$141
Xnfet$162_15 m1_14556_21786# m1_14556_21786# vss vss m1_13394_21586# vss nfet$162
Xpfet$145_10 vdd vdd m1_27031_17343# m1_n10452_25858# pfet$145
Xpfet$166_9 vdd vdd m1_n4464_25980# m1_n4623_25487# pfet$166
Xnfet$154_16 m1_26873_21786# vss m1_27003_21590# vss nfet$154
Xnfet$170_15 m1_17697_15478# m1_17697_15478# m1_n2543_20130# m1_n2543_20130# m1_20407_20470#
+ vss nfet$170
Xnfet$172_5 m1_27031_17343# m1_29087_15778# m1_28470_16080# vss nfet$172
Xnfet$158_3 m1_n7513_20152# vss m1_326_24346# vss nfet$158
Xpfet$142_33 vdd m1_28490_22513# m1_28490_22513# m1_27462_22102# m1_29256_21786# m1_29256_21786#
+ pfet$142
Xpfet$142_22 vdd m1_21456_22513# m1_21456_22513# m1_20428_22102# m1_22222_21786# m1_22222_21786#
+ pfet$142
Xpfet$164_6 vdd m1_n10308_24542# vdd m1_n9336_24346# pfet$164
Xpfet$142_11 vdd vdd vdd m1_2843_22102# m1_2384_21590# m1_2384_21590# pfet$142
Xnfet$149_27 m1_12875_24346# m1_12875_24346# vss vss m1_12357_24542# vss nfet$149
Xnfet$149_16 m1_24808_24224# m1_24808_24224# m1_24452_24542# m1_24452_24542# m1_24906_24542#
+ vss nfet$149
Xnfet$163_1 m1_14422_22513# m1_14422_22513# m1_31535_19792# m1_31535_19792# m1_31771_20470#
+ vss nfet$163
Xnfet$170_2 m1_n3218_15478# m1_n3218_15478# m1_2590_19404# m1_2590_19404# m1_2822_20470#
+ vss nfet$170
Xnfet$156_0 sd9 vss m1_n7401_15478# vss nfet$156
Xpfet$162_3 vdd m1_n3184_24224# m1_n3651_26174# m1_n4623_25487# pfet$162
Xnfet$151_17 m1_12935_21590# m1_12935_21590# m1_14422_22513# m1_14422_22513# m1_13394_21586#
+ vss nfet$151
Xpfet$148_1 vdd vdd m1_n1134_25662# m1_n1271_25858# pfet$148
Xpfet$141_8 vdd vdd m1_9331_15478# sd5 pfet$141
Xpfet$148_10 vdd vdd m1_35071_24542# m1_32675_25947# pfet$148
Xpfet$160_0 vdd vdd m1_n7513_20152# m1_35837_22102# pfet$160
Xnfet$162_16 m1_28624_21786# m1_28624_21786# vss vss m1_27462_21586# vss nfet$162
Xpfet$145_11 vdd vdd m1_26807_17518# m1_26217_17714# pfet$145
Xnfet$154_17 m1_25107_21786# vss m1_25739_21786# vss nfet$154
Xnfet$170_16 m1_25722_20152# m1_25722_20152# m1_n3206_20274# m1_n3206_20274# m1_24556_20470#
+ vss nfet$170
Xnfet$172_6 m1_27190_17836# m1_28113_15778# m1_27292_16202# vss nfet$172
Xnfet$158_4 m1_n789_25858# vss m1_1607_24542# vss nfet$158
Xpfet$142_34 vdd vdd vdd m1_28090_22402# m1_26873_21786# m1_26873_21786# pfet$142
Xpfet$142_23 vdd vdd vdd m1_23945_22102# m1_23486_21590# m1_23486_21590# pfet$142
Xpfet$164_7 vdd vdd m1_n10452_25858# m1_n4978_24224# pfet$164
Xpfet$142_12 vdd vdd vdd m1_3471_22402# m1_2254_21786# m1_2254_21786# pfet$142
Xnfet$149_17 m1_20625_24224# m1_20625_24224# m1_20269_24542# m1_20269_24542# m1_20723_24542#
+ vss nfet$149
Xnfet$156_1 sd2 vss m1_21880_15478# vss nfet$156
Xnfet$163_2 m1_17939_22513# m1_17939_22513# vss vss m1_31771_20470# vss nfet$163
Xnfet$170_3 m1_8137_20152# m1_8137_20152# m1_6107_19404# m1_6107_19404# m1_6971_20470#
+ vss nfet$170
Xnfet$149_0 m1_4509_24346# m1_4509_24346# vss vss m1_3991_24542# vss nfet$149
Xpfet$162_4 vdd m1_n2567_23922# m1_n3184_24224# m1_n4464_25980# pfet$162
Xpfet$148_2 vdd vdd m1_n1271_25858# m1_n10452_25858# pfet$148
Xpfet$141_9 vdd vdd m1_8172_15778# m1_5302_17714# pfet$141
Xpfet$148_11 vdd vdd m1_32817_25662# m1_32675_25947# pfet$148
Xpfet$153_0 vdd vdd m1_n1263_21786# pd1 pfet$153
Xnfet$162_17 m1_29256_21786# m1_29256_21786# vss vss m1_28094_21586# vss nfet$162
Xpfet$145_12 vdd vdd m1_26676_16080# m1_n7513_20152# pfet$145
Xnfet$179_0 m1_n10933_25858# m1_n8848_25658# m1_n8055_24542# vss nfet$179
Xnfet$170_17 m1_21880_15478# m1_21880_15478# m1_n3206_20274# m1_n3206_20274# m1_23924_20470#
+ vss nfet$170
Xnfet$172_7 m1_27190_17836# m1_28470_16080# m1_28003_18030# vss nfet$172
Xnfet$158_5 m1_n789_25858# vss m1_488_21786# vss nfet$158
Xpfet$142_35 vdd vdd vdd m1_13394_22102# m1_12935_21590# m1_12935_21590# pfet$142
Xnfet$149_18 m1_21241_24346# m1_21241_24346# vss vss m1_20723_24542# vss nfet$149
Xpfet$142_24 vdd m1_17939_22513# m1_17939_22513# m1_16911_22102# m1_18705_21786# m1_18705_21786#
+ pfet$142
Xpfet$142_13 vdd vdd vdd m1_6988_22402# m1_5771_21786# m1_5771_21786# pfet$142
Xnfet$156_2 sd1 vss m1_26063_15478# vss nfet$156
Xnfet$163_3 m1_24973_22513# m1_24973_22513# vss vss m1_30492_20470# vss nfet$163
Xnfet$170_4 m1_965_15478# m1_965_15478# m1_6107_19404# m1_6107_19404# m1_6339_20470#
+ vss nfet$170
Xnfet$149_1 m1_3893_24224# m1_3893_24224# m1_3537_24542# m1_3537_24542# m1_3991_24542#
+ vss nfet$149
Xpfet$148_3 vdd vdd m1_1607_24542# m1_n789_25858# pfet$148
Xpfet$162_5 vdd m1_n10572_23922# m1_n10308_24542# m1_n10933_25858# pfet$162
Xpfet$148_12 vdd vdd m1_32193_25858# m1_25107_21786# pfet$148
Xnfet$161_0 m1_n290_24224# m1_n290_24224# m1_n646_24542# m1_n646_24542# m1_n192_24542#
+ vss nfet$161
Xpfet$153_1 vdd vdd m1_2254_21786# pd2 pfet$153
Xpfet$146_0 vdd vdd m1_2384_19550# m1_n3534_17714# pfet$146
Xpfet$140_90 vdd vdd m1_24309_25858# m1_25424_24346# pfet$140
Xpfet$145_13 vdd vdd m1_25747_17714# m1_26217_17714# pfet$145
Xnfet$179_1 m1_n10796_25662# m1_n10572_23922# m1_n10308_24542# vss nfet$179
Xnfet$158_6 m1_n910_23922# vss m1_n290_24224# vss nfet$158
Xnfet$149_19 m1_21729_25658# m1_21729_25658# vss vss m1_22188_25502# vss nfet$149
Xpfet$142_25 vdd m1_17939_22513# m1_17939_22513# m1_17539_22402# m1_18073_21786# m1_18073_21786#
+ pfet$142
Xpfet$142_14 vdd vdd vdd m1_n46_22402# m1_n1263_21786# m1_n1263_21786# pfet$142
Xnfet$163_4 m1_32818_20470# m1_32818_20470# vss vss m1_34329_20470# vss nfet$163
Xnfet$149_2 m1_4997_25658# m1_4997_25658# vss vss m1_5456_25502# vss nfet$149
Xnfet$170_5 m1_5148_15478# m1_5148_15478# m1_9624_19404# m1_9624_19404# m1_9856_20470#
+ vss nfet$170
Xpfet$148_4 vdd vdd m1_488_21786# m1_n789_25858# pfet$148
Xpfet$162_6 vdd m1_n8848_25658# m1_n8055_24542# m1_n10796_25662# pfet$162
Xnfet$161_1 m1_814_25658# m1_814_25658# vss vss m1_1273_25502# vss nfet$161
Xnfet$154_0 m1_n1263_21786# vss m1_n1133_21590# vss nfet$154
Xpfet$148_13 vdd vdd m1_33790_24346# m1_n7513_20152# pfet$148
Xpfet$153_2 vdd vdd m1_26873_21786# pd9 pfet$153
Xpfet$146_1 vdd vdd m1_4620_20152# m1_n3218_15478# pfet$146
Xpfet$140_91 vdd vdd m1_23356_21786# pd8 pfet$140
Xpfet$140_80 vdd vdd m1_17058_24346# m1_n7513_20152# pfet$140
Xnfet$179_2 m1_n10933_25858# m1_n10309_25662# m1_n10572_23922# vss nfet$179
Xnfet$158_7 m1_25107_21786# vss m1_32193_25858# vss nfet$158
Xpfet$142_26 vdd vdd vdd m1_16911_22102# m1_16452_21590# m1_16452_21590# pfet$142
Xpfet$142_15 vdd m1_354_22513# m1_354_22513# m1_n46_22402# m1_488_21786# m1_488_21786#
+ pfet$142
Xnfet$184_0 m1_n4485_20152# m1_n6380_21786# vss vss nfet$184
Xpfet$169_0 vdd m1_n6380_21786# m1_n6380_21786# m1_n5019_19550# m1_n5227_20152# m1_n5227_20152#
+ pfet$169
Xnfet$170_6 m1_11654_20152# m1_11654_20152# m1_9624_19404# m1_9624_19404# m1_10488_20470#
+ vss nfet$170
Xnfet$163_5 m1_32818_21586# m1_32818_21586# m1_34093_19792# m1_34093_19792# m1_34329_20470#
+ vss nfet$163
Xpfet$148_5 vdd vdd m1_326_24346# m1_n7513_20152# pfet$148
Xnfet$149_3 m1_4509_24346# m1_4509_24346# m1_3394_25858# m1_3394_25858# m1_5456_25502#
+ vss nfet$149
Xpfet$162_7 vdd m1_n3541_23922# m1_n4362_24346# m1_n4623_25487# pfet$162
Xnfet$161_2 m1_326_24346# m1_326_24346# m1_n789_25858# m1_n789_25858# m1_1273_25502#
+ vss nfet$161
Xnfet$154_1 m1_11039_21786# vss m1_11671_21786# vss nfet$154
Xpfet$146_2 vdd vdd m1_1103_20152# m1_n7401_15478# pfet$146
Xpfet$140_92 vdd vdd m1_28492_25858# m1_29607_24346# pfet$140
Xpfet$140_81 vdd vdd m1_18339_24542# m1_15943_25858# pfet$140
Xpfet$140_70 vdd vdd m1_14156_24542# m1_11760_25858# pfet$140
Xpfet$151_0 vdd m1_31535_19792# vdd m1_17939_22513# pfet$151
Xnfet$179_3 m1_n10796_25662# m1_n9952_24224# m1_n8848_25658# vss nfet$179
Xnfet$158_8 m1_32193_25858# vss m1_32330_25662# vss nfet$158
Xpfet$142_27 vdd m1_14422_22513# m1_14422_22513# m1_14022_22402# m1_14556_21786# m1_14556_21786#
+ pfet$142
Xpfet$142_16 vdd m1_24973_22513# m1_24973_22513# m1_23945_22102# m1_25739_21786# m1_25739_21786#
+ pfet$142
Xnfet$184_1 m1_n5227_20152# vss m1_n6380_21786# vss nfet$184
Xnfet$177_0 m1_n8625_26174# vss m1_n8055_24542# vss nfet$177
Xpfet$169_1 vdd vdd vdd m1_n5019_22344# m1_n4485_21904# m1_n4485_21904# pfet$169
Xnfet$163_6 m1_354_22513# m1_354_22513# m1_31535_22102# m1_31535_22102# m1_31771_21430#
+ vss nfet$163
Xnfet$170_7 m1_n7401_15478# m1_n7401_15478# m1_n927_19404# m1_n927_19404# m1_n695_20470#
+ vss nfet$170
Xnfet$149_4 m1_12259_24224# m1_12259_24224# m1_11903_24542# m1_11903_24542# m1_12357_24542#
+ vss nfet$149
Xpfet$148_6 vdd vdd m1_n290_24224# m1_n910_23922# pfet$148
Xnfet$161_3 m1_326_24346# m1_326_24346# vss vss m1_n192_24542# vss nfet$161
Xnfet$154_2 m1_12805_21786# vss m1_12935_21590# vss nfet$154
Xpfet$146_3 vdd vdd m1_5901_19550# m1_649_17714# pfet$146
Xnfet$152_10 m1_9015_17714# m1_9015_17714# vss vss m1_14005_20470# vss nfet$152
Xpfet$140_93 vdd m1_28991_24224# m1_30095_25658# m1_28010_25858# pfet$140
Xpfet$140_82 vdd vdd m1_21241_24346# m1_n7513_20152# pfet$140
Xpfet$140_71 vdd vdd m1_11039_21786# m1_11760_25858# pfet$140
Xpfet$140_60 vdd vdd m1_20126_25858# m1_21241_24346# pfet$140
Xpfet$151_1 vdd vdd m1_30256_19792# m1_21456_22513# pfet$151
Xpfet$144_0 vdd vdd m1_n1133_21590# m1_n1263_21786# pfet$144
Xnfet$179_4 m1_n4623_25487# m1_n2567_23922# m1_n3184_24224# vss nfet$179
Xnfet$158_9 m1_n7513_20152# vss m1_33790_24346# vss nfet$158
Xpfet$142_28 vdd m1_14422_22513# m1_14422_22513# m1_13394_22102# m1_15188_21786# m1_15188_21786#
+ pfet$142
Xpfet$142_17 vdd m1_21456_22513# m1_21456_22513# m1_21056_22402# m1_21590_21786# m1_21590_21786#
+ pfet$142
Xnfet$177_1 m1_n8625_26174# vss m1_n7082_23622# vss nfet$177
Xpfet$169_2 vdd m1_n5764_21786# m1_n5764_21786# m1_n5019_22344# m1_n5227_21418# m1_n5227_21418#
+ pfet$169
Xnfet$163_7 m1_3871_22513# m1_3871_22513# vss vss m1_31771_21430# vss nfet$163
Xnfet$155_10 m1_26063_15478# vss m1_29239_20152# vss nfet$155
Xnfet$170_8 m1_26063_15478# m1_26063_15478# m1_n3822_20130# m1_n3822_20130# m1_27441_20470#
+ vss nfet$170
Xnfet$149_5 m1_8692_24346# m1_8692_24346# vss vss m1_8174_24542# vss nfet$149
Xpfet$148_7 vdd vdd m1_32330_25662# m1_32193_25858# pfet$148
Xnfet$161_4 m1_33174_24224# m1_33174_24224# m1_32818_24542# m1_32818_24542# m1_33272_24542#
+ vss nfet$161
Xpfet$146_4 vdd vdd m1_12935_19550# m1_9015_17714# pfet$146
Xnfet$154_3 m1_9288_21786# vss m1_9418_21590# vss nfet$154
Xnfet$152_11 m1_13198_17714# m1_13198_17714# vss vss m1_17522_20470# vss nfet$152
Xnfet$152_0 m1_n3534_17714# m1_n3534_17714# vss vss m1_3454_20470# vss nfet$152
Xpfet$151_2 vdd m1_30256_19792# vdd m1_24973_22513# pfet$151
Xpfet$144_1 vdd vdd m1_11671_21786# m1_11039_21786# pfet$144
Xpfet$140_94 vdd m1_28492_25858# vdd m1_30095_25658# pfet$140
Xpfet$140_83 vdd m1_21729_25658# m1_22522_24542# m1_19781_25662# pfet$140
Xpfet$140_72 vdd m1_13363_25658# m1_14156_24542# m1_11415_25662# pfet$140
Xpfet$140_61 vdd m1_24452_24542# vdd m1_25424_24346# pfet$140
Xpfet$140_50 vdd vdd m1_20268_25662# m1_20126_25858# pfet$140
Xnfet$158_10 m1_32675_25947# vss m1_35071_24542# vss nfet$158
Xnfet$179_5 m1_n4464_25980# m1_n3541_23922# m1_n4362_24346# vss nfet$179
Xnfet$169_20 m1_22493_16080# m1_22493_16080# m1_22034_17714# m1_22034_17714# m1_22591_16398#
+ vss nfet$169
Xnfet$177_2 vss vss m1_n9336_24346# vss nfet$177
Xpfet$142_29 vdd vdd vdd m1_14022_22402# m1_12805_21786# m1_12805_21786# pfet$142
Xpfet$142_18 vdd vdd vdd m1_24573_22402# m1_23356_21786# m1_23356_21786# pfet$142
Xnfet$155_11 m1_9331_15478# vss m1_15171_20152# vss nfet$155
Xnfet$170_9 m1_29239_20152# m1_29239_20152# m1_n3822_20130# m1_n3822_20130# m1_28073_20470#
+ vss nfet$170
Xnfet$149_6 m1_8076_24224# m1_8076_24224# m1_7720_24542# m1_7720_24542# m1_8174_24542#
+ vss nfet$149
Xpfet$148_8 vdd vdd m1_33174_24224# m1_32554_23922# pfet$148
Xnfet$182_0 m1_n4485_21904# m1_n5764_21786# vss vss nfet$182
Xpfet$167_0 vdd vdd m1_n7186_25858# m1_n10452_25858# pfet$167
Xnfet$161_5 m1_33790_24346# m1_33790_24346# vss vss m1_33272_24542# vss nfet$161
Xnfet$154_4 m1_7522_21786# vss m1_8154_21786# vss nfet$154
Xpfet$146_5 vdd vdd m1_8137_20152# m1_965_15478# pfet$146
Xnfet$152_12 m1_16452_19550# m1_16452_19550# vss vss m1_16890_20470# vss nfet$152
Xpfet$151_3 vdd vdd m1_34843_21786# m1_34093_19792# pfet$151
Xnfet$152_1 m1_2384_19550# m1_2384_19550# vss vss m1_2822_20470# vss nfet$152
Xpfet$144_2 vdd vdd m1_12935_21590# m1_12805_21786# pfet$144
Xpfet$140_95 vdd vdd m1_28991_24224# m1_28371_23922# pfet$140
Xpfet$140_84 vdd vdd m1_23827_25858# m1_18073_21786# pfet$140
Xpfet$140_73 vdd m1_16086_24542# vdd m1_17058_24346# pfet$140
Xpfet$140_62 vdd vdd m1_24452_24542# m1_24808_24224# pfet$140
Xpfet$140_51 vdd vdd m1_20625_24224# m1_20005_23922# pfet$140
Xpfet$140_40 vdd vdd m1_11760_25858# m1_12875_24346# pfet$140
Xnfet$158_11 m1_32554_23922# vss m1_33174_24224# vss nfet$158
Xnfet$179_6 m1_n4464_25980# m1_n3184_24224# m1_n3651_26174# vss nfet$179
Xnfet$169_10 m1_1578_16080# m1_1578_16080# m1_1119_17714# m1_1119_17714# m1_1676_16398#
+ vss nfet$169
Xnfet$177_3 fin vss m1_n10933_25858# vss nfet$177
Xpfet$142_19 vdd m1_24973_22513# m1_24973_22513# m1_24573_22402# m1_25107_21786# m1_25107_21786#
+ pfet$142
Xnfet$169_21 m1_14127_16080# m1_14127_16080# vss vss m1_15690_17358# vss nfet$169
Xnfet$149_7 m1_9180_25658# m1_9180_25658# vss vss m1_9639_25502# vss nfet$149
Xpfet$148_9 vdd vdd m1_28624_21786# m1_32675_25947# pfet$148
Xnfet$155_12 m1_13514_15478# vss m1_18688_20152# vss nfet$155
Xnfet$182_1 m1_n5227_21418# vss m1_n5764_21786# vss nfet$182
Xnfet$175_0 m1_n7082_23622# m1_n6856_24542# vss vss nfet$175
Xpfet$167_1 vdd m1_n7186_25858# vdd m1_n6111_25858# pfet$167
Xnfet$161_6 m1_33790_24346# m1_33790_24346# m1_32675_25947# m1_32675_25947# m1_34737_25502#
+ vss nfet$161
Xnfet$154_5 m1_488_21786# vss m1_1120_21786# vss nfet$154
Xpfet$146_6 vdd vdd m1_9418_19550# m1_4832_17714# pfet$146
Xnfet$152_13 m1_19969_19550# m1_19969_19550# vss vss m1_20407_20470# vss nfet$152
Xpfet$151_4 vdd m1_34093_19792# vdd m1_32818_20470# pfet$151
Xnfet$152_2 m1_5901_19550# m1_5901_19550# vss vss m1_6339_20470# vss nfet$152
Xnfet$177_10 vss vss m1_n4978_24224# vss nfet$177
Xpfet$144_3 vdd vdd m1_9418_21590# m1_9288_21786# pfet$144
Xpfet$140_96 vdd m1_28635_24542# vdd m1_29607_24346# pfet$140
Xpfet$140_85 vdd m1_24188_23922# m1_24452_24542# m1_23827_25858# pfet$140
Xpfet$140_74 vdd vdd m1_14556_21786# m1_15943_25858# pfet$140
Xpfet$140_63 vdd vdd m1_19781_25662# m1_19644_25858# pfet$140
Xpfet$140_52 vdd m1_20268_25662# m1_20005_23922# m1_19781_25662# pfet$140
Xpfet$140_41 vdd vdd m1_9288_21786# pd4 pfet$140
Xpfet$140_30 vdd vdd m1_2912_25858# m1_488_21786# pfet$140
Xpfet$142_0 vdd vdd vdd m1_n674_22102# m1_n1133_21590# m1_n1133_21590# pfet$142
Xnfet$158_12 m1_32675_25947# vss m1_28624_21786# vss nfet$158
Xnfet$179_7 m1_n4623_25487# m1_n4362_24346# m1_n4847_25662# vss nfet$179
Xpfet$141_110 vdd vdd m1_10458_17836# m1_10299_17343# pfet$141
Xnfet$169_22 m1_15564_15778# m1_15564_15778# m1_15454_18030# m1_15454_18030# m1_15690_17358#
+ vss nfet$169
Xnfet$169_11 m1_6377_16202# m1_6377_16202# vss vss m1_5859_16398# vss nfet$169
Xnfet$177_4 m1_n10572_23922# vss m1_n9952_24224# vss nfet$177
Xnfet$168_0 fout vss m1_35837_22102# vss nfet$168
Xnfet$155_13 m1_13198_17714# vss m1_16452_19550# vss nfet$155
Xnfet$149_8 m1_8692_24346# m1_8692_24346# m1_7577_25858# m1_7577_25858# m1_9639_25502#
+ vss nfet$149
Xnfet$182_2 m1_n6839_21786# vss m1_n6973_21481# vss nfet$182
Xnfet$175_1 m1_n8283_19850# vss m1_n6856_24542# vss nfet$175
Xpfet$143_30 vdd vdd vdd m1_24560_19550# m1_21880_15478# m1_21880_15478# pfet$143
Xnfet$161_7 m1_34278_25658# m1_34278_25658# vss vss m1_34737_25502# vss nfet$161
Xnfet$154_6 m1_5771_21786# vss m1_5901_21590# vss nfet$154
Xpfet$146_7 vdd vdd m1_11654_20152# m1_5148_15478# pfet$146
Xnfet$152_14 m1_17381_17714# m1_17381_17714# vss vss m1_21039_20470# vss nfet$152
Xpfet$172_0 vdd vdd m1_n8145_21908# m1_n6839_20152# pfet$172
Xnfet$152_3 m1_4832_17714# m1_4832_17714# vss vss m1_10488_20470# vss nfet$152
Xnfet$177_11 m1_n10452_25858# vss m1_n4847_25662# vss nfet$177
Xpfet$140_97 vdd vdd m1_21590_21786# m1_24309_25858# pfet$140
Xpfet$140_86 vdd m1_28634_25662# m1_28371_23922# m1_28147_25662# pfet$140
Xpfet$140_75 vdd vdd m1_19644_25858# m1_14556_21786# pfet$140
Xpfet$140_64 vdd vdd m1_22522_24542# m1_20126_25858# pfet$140
Xpfet$140_53 vdd m1_20625_24224# m1_21729_25658# m1_19644_25858# pfet$140
Xpfet$140_42 vdd m1_11760_25858# vdd m1_13363_25658# pfet$140
Xpfet$151_5 vdd vdd m1_34093_19792# m1_32818_21586# pfet$151
Xpfet$140_31 vdd m1_3273_23922# m1_3537_24542# m1_2912_25858# pfet$140
Xpfet$140_20 vdd vdd m1_4509_24346# m1_n7513_20152# pfet$140
Xpfet$144_4 vdd vdd m1_8154_21786# m1_7522_21786# pfet$144
Xpfet$142_1 vdd m1_7388_22513# m1_7388_22513# m1_6988_22402# m1_7522_21786# m1_7522_21786#
+ pfet$142
Xnfet$150_0 m1_3394_25858# vss m1_5790_24542# vss nfet$150
Xnfet$158_13 m1_32675_25947# vss m1_32817_25662# vss nfet$158
Xpfet$141_100 vdd vdd m1_23820_18030# m1_23930_15778# pfet$141
Xnfet$169_23 m1_18926_16202# m1_18926_16202# vss vss m1_18408_16398# vss nfet$169
Xnfet$169_12 m1_n1168_15778# m1_n1168_15778# m1_n1278_18030# m1_n1278_18030# m1_n1042_17358#
+ vss nfet$169
Xnfet$177_5 m1_n10933_25858# vss m1_n10796_25662# vss nfet$177
Xnfet$150_80 m1_28147_25662# m1_28991_24224# m1_30095_25658# vss nfet$150
Xnfet$149_9 m1_17058_24346# m1_17058_24346# vss vss m1_16540_24542# vss nfet$149
Xnfet$155_14 m1_21564_17714# vss m1_23486_19550# vss nfet$155
Xnfet$168_1 define m1_35837_22102# vss vss nfet$168
Xpfet$143_31 vdd m1_n2543_20130# m1_n2543_20130# m1_20407_19850# m1_19969_19550# m1_19969_19550#
+ pfet$143
Xpfet$143_20 vdd m1_n3822_21786# m1_n3822_21786# m1_14009_19550# m1_9015_17714# m1_9015_17714#
+ pfet$143
Xnfet$154_7 m1_4005_21786# vss m1_4637_21786# vss nfet$154
Xpfet$146_8 vdd vdd m1_n1133_19550# m1_n7383_17599# pfet$146
Xnfet$180_0 m1_n7186_25858# vss m1_n7320_25516# vss nfet$180
Xpfet$165_0 vdd vdd m1_n4485_20152# m1_n3822_20130# pfet$165
Xnfet$152_15 m1_21564_17714# m1_21564_17714# vss vss m1_24556_20470# vss nfet$152
Xnfet$152_4 m1_9418_19550# m1_9418_19550# vss vss m1_9856_20470# vss nfet$152
Xnfet$177_12 m1_n10452_25858# vss m1_n5571_25662# vss nfet$177
Xpfet$140_98 vdd m1_30095_25658# m1_30888_24542# m1_28147_25662# pfet$140
Xpfet$140_87 vdd vdd m1_28147_25662# m1_28010_25858# pfet$140
Xpfet$140_76 vdd m1_20005_23922# m1_20269_24542# m1_19644_25858# pfet$140
Xpfet$140_65 vdd vdd m1_18073_21786# m1_20126_25858# pfet$140
Xpfet$140_54 vdd vdd m1_24808_24224# m1_24188_23922# pfet$140
Xpfet$140_43 vdd vdd m1_12805_21786# pd5 pfet$140
Xpfet$151_6 vdd vdd m1_31535_19792# m1_14422_22513# pfet$151
Xpfet$140_32 vdd vdd m1_7720_24542# m1_8076_24224# pfet$140
Xpfet$140_21 vdd m1_7456_23922# m1_7720_24542# m1_7095_25858# pfet$140
Xpfet$140_10 vdd m1_8076_24224# m1_9180_25658# m1_7095_25858# pfet$140
Xpfet$144_5 vdd vdd m1_1120_21786# m1_488_21786# pfet$144
Xnfet$153_80 m1_18824_17836# m1_19747_15778# m1_18926_16202# vss nfet$153
Xpfet$142_2 vdd m1_7388_22513# m1_7388_22513# m1_6360_22102# m1_8154_21786# m1_8154_21786#
+ pfet$142
Xnfet$150_1 m1_2912_25858# m1_4997_25658# m1_5790_24542# vss nfet$150
Xpfet$141_101 vdd vdd m1_19637_18030# m1_19747_15778# pfet$141
Xnfet$169_24 m1_18310_16080# m1_18310_16080# m1_17851_17714# m1_17851_17714# m1_18408_16398#
+ vss nfet$169
Xnfet$169_13 m1_n2605_16080# m1_n2605_16080# vss vss m1_n1042_17358# vss nfet$169
Xnfet$177_6 m1_n10452_25858# vss m1_n10309_25662# vss nfet$177
Xnfet$150_81 m1_n7513_20152# vss m1_25424_24346# vss nfet$150
Xnfet$150_70 m1_21590_21786# vss m1_28010_25858# vss nfet$150
Xnfet$155_15 m1_17697_15478# vss m1_22205_20152# vss nfet$155
Xpfet$143_32 vdd m1_n2543_20130# m1_n2543_20130# m1_21043_19550# m1_17381_17714# m1_17381_17714#
+ pfet$143
Xpfet$143_21 vdd vdd vdd m1_13373_19850# m1_15171_20152# m1_15171_20152# pfet$143
Xpfet$143_10 vdd vdd vdd m1_9856_19850# m1_11654_20152# m1_11654_20152# pfet$143
Xpfet$146_9 vdd vdd m1_27003_19550# m1_25747_17714# pfet$146
Xnfet$173_0 m1_n5351_15778# m1_n5351_15778# m1_n5461_18030# m1_n5461_18030# m1_n5225_17358#
+ vss nfet$173
Xnfet$180_1 m1_n6856_24542# vss m1_n6111_25858# vss nfet$180
Xnfet$154_8 m1_2254_21786# vss m1_2384_21590# vss nfet$154
Xpfet$158_0 vdd vdd m1_n7247_17714# m1_n6788_16080# pfet$158
Xpfet$165_1 vdd m1_n4485_21904# vdd m1_9624_19404# pfet$165
Xnfet$152_16 m1_23486_19550# m1_23486_19550# vss vss m1_23924_20470# vss nfet$152
Xnfet$152_5 m1_649_17714# m1_649_17714# vss vss m1_6971_20470# vss nfet$152
Xnfet$177_13 fin vss m1_n4623_25487# vss nfet$177
Xpfet$151_7 vdd vdd m1_31535_22102# m1_354_22513# pfet$151
Xpfet$140_33 vdd vdd m1_7522_21786# m1_7577_25858# pfet$140
Xpfet$140_22 vdd vdd m1_3537_24542# m1_3893_24224# pfet$140
Xpfet$140_11 vdd vdd m1_7719_25662# m1_7577_25858# pfet$140
Xpfet$144_6 vdd vdd m1_5901_21590# m1_5771_21786# pfet$144
Xpfet$140_99 vdd vdd m1_26705_24542# m1_24309_25858# pfet$140
Xpfet$140_88 vdd vdd m1_28634_25662# m1_28492_25858# pfet$140
Xpfet$140_77 vdd vdd m1_20269_24542# m1_20625_24224# pfet$140
Xpfet$140_66 vdd vdd m1_15461_25858# m1_11039_21786# pfet$140
Xpfet$140_55 vdd m1_24451_25662# m1_24188_23922# m1_23964_25662# pfet$140
Xpfet$140_44 vdd m1_15943_25858# vdd m1_17546_25658# pfet$140
Xnfet$153_81 m1_13198_17714# vss m1_10299_17343# vss nfet$153
Xnfet$153_70 m1_n7513_20152# vss m1_18310_16080# vss nfet$153
Xnfet$150_2 m1_n7513_20152# vss m1_4509_24346# vss nfet$150
Xpfet$142_3 vdd m1_9645_21447# m1_9645_21447# m1_10505_22402# m1_11039_21786# m1_11039_21786#
+ pfet$142
Xpfet$146_10 vdd vdd m1_29239_20152# m1_26063_15478# pfet$146
Xpfet$140_0 vdd vdd m1_3049_25662# m1_2912_25858# pfet$140
Xpfet$141_102 vdd vdd m1_13198_17714# m1_13668_17714# pfet$141
Xnfet$169_25 m1_14743_16202# m1_14743_16202# vss vss m1_14225_16398# vss nfet$169
Xnfet$169_14 m1_n2605_16080# m1_n2605_16080# m1_n3064_17714# m1_n3064_17714# m1_n2507_16398#
+ vss nfet$169
Xnfet$177_7 m1_n7320_25516# vss m1_n2567_23922# vss nfet$177
Xnfet$150_82 m1_11415_25662# m1_12259_24224# m1_13363_25658# vss nfet$150
Xnfet$150_71 m1_28147_25662# m1_28371_23922# m1_28635_24542# vss nfet$150
Xnfet$150_60 pd6 vss m1_16322_21786# vss nfet$150
Xnfet$155_16 m1_17381_17714# vss m1_19969_19550# vss nfet$155
Xpfet$143_33 vdd m1_n3206_20274# m1_n3206_20274# m1_24560_19550# m1_21564_17714# m1_21564_17714#
+ pfet$143
Xpfet$143_22 vdd vdd vdd m1_14009_19550# m1_9331_15478# m1_9331_15478# pfet$143
Xpfet$143_11 vdd vdd vdd m1_10492_19550# m1_5148_15478# m1_5148_15478# pfet$143
Xnfet$154_9 m1_23356_21786# vss m1_23486_21590# vss nfet$154
Xnfet$166_0 m1_34093_19792# vss m1_34843_21786# vss nfet$166
Xnfet$173_1 m1_n6788_16080# m1_n6788_16080# vss vss m1_n5225_17358# vss nfet$173
Xpfet$158_1 vdd m1_n7247_17714# vdd m1_n6172_16202# pfet$158
Xpfet$165_2 vdd m1_n5227_21418# vdd m1_2590_19404# pfet$165
Xnfet$152_17 m1_12935_19550# m1_12935_19550# vss vss m1_13373_20470# vss nfet$152
Xnfet$152_6 m1_n1133_19550# m1_n1133_19550# vss vss m1_n695_20470# vss nfet$152
Xpfet$144_7 vdd vdd m1_4637_21786# m1_4005_21786# pfet$144
Xpfet$140_89 vdd vdd m1_19839_21786# pd7 pfet$140
Xpfet$140_78 vdd m1_20269_24542# vdd m1_21241_24346# pfet$140
Xpfet$140_67 vdd m1_15822_23922# m1_16086_24542# m1_15461_25858# pfet$140
Xpfet$140_56 vdd m1_24808_24224# m1_25912_25658# m1_23827_25858# pfet$140
Xpfet$140_45 vdd vdd m1_16442_24224# m1_15822_23922# pfet$140
Xpfet$140_34 vdd m1_9180_25658# m1_9973_24542# m1_7232_25662# pfet$140
Xpfet$140_23 vdd m1_3537_24542# vdd m1_4509_24346# pfet$140
Xpfet$140_12 vdd m1_7577_25858# vdd m1_9180_25658# pfet$140
Xpfet$170_0 vdd vdd m1_n5227_20152# m1_n2543_20130# pfet$170
Xnfet$150_3 m1_488_21786# vss m1_2912_25858# vss nfet$150
Xnfet$153_82 m1_10299_17343# vss m1_10458_17836# vss nfet$153
Xnfet$153_71 m1_14641_17836# m1_15921_16080# m1_15454_18030# vss nfet$153
Xnfet$153_60 m1_18665_17343# vss m1_18824_17836# vss nfet$153
Xpfet$142_4 vdd vdd vdd m1_9877_22102# m1_9418_21590# m1_9418_21590# pfet$142
Xpfet$141_103 vdd m1_14743_16202# m1_14258_17518# m1_14641_17836# pfet$141
Xpfet$146_11 vdd vdd m1_18688_20152# m1_13514_15478# pfet$146
Xnfet$169_26 m1_14127_16080# m1_14127_16080# m1_13668_17714# m1_13668_17714# m1_14225_16398#
+ vss nfet$169
Xpfet$140_1 vdd m1_3536_25662# m1_3273_23922# m1_3049_25662# pfet$140
Xnfet$169_15 m1_n1989_16202# m1_n1989_16202# vss vss m1_n2507_16398# vss nfet$169
Xnfet$177_8 m1_n4623_25487# vss m1_n4464_25980# vss nfet$177
Xnfet$150_72 m1_23827_25858# m1_25912_25658# m1_26705_24542# vss nfet$150
Xnfet$150_61 m1_23964_25662# m1_24808_24224# m1_25912_25658# vss nfet$150
Xnfet$150_50 m1_n7513_20152# vss m1_21241_24346# vss nfet$150
Xnfet$155_17 m1_21880_15478# vss m1_25722_20152# vss nfet$155
Xpfet$143_34 vdd m1_n3206_20274# m1_n3206_20274# m1_23924_19850# m1_23486_19550# m1_23486_19550#
+ pfet$143
Xpfet$143_23 vdd vdd vdd m1_16890_19850# m1_18688_20152# m1_18688_20152# pfet$143
Xpfet$143_12 vdd m1_6107_19404# m1_6107_19404# m1_6975_19550# m1_649_17714# m1_649_17714#
+ pfet$143
Xnfet$166_1 m1_30256_19792# vss m1_32818_20470# vss nfet$166
Xnfet$173_2 m1_n6788_16080# m1_n6788_16080# m1_n7247_17714# m1_n7247_17714# m1_n6690_16398#
+ vss nfet$173
Xpfet$165_3 vdd vdd m1_n5227_21418# m1_6107_19404# pfet$165
Xnfet$159_0 m1_n1134_25662# m1_n910_23922# m1_n646_24542# vss nfet$159
Xpfet$158_2 vdd vdd m1_n5461_18030# m1_n5351_15778# pfet$158
Xnfet$152_7 m1_n7383_17599# m1_n7383_17599# vss vss m1_n63_20470# vss nfet$152
Xpfet$144_8 vdd vdd m1_2384_21590# m1_2254_21786# pfet$144
Xpfet$140_79 vdd m1_17546_25658# m1_18339_24542# m1_15598_25662# pfet$140
Xpfet$140_68 vdd vdd m1_16086_24542# m1_16442_24224# pfet$140
Xpfet$140_57 vdd vdd m1_24451_25662# m1_24309_25858# pfet$140
Xpfet$140_46 vdd m1_16442_24224# m1_17546_25658# m1_15461_25858# pfet$140
Xpfet$140_35 vdd m1_7720_24542# vdd m1_8692_24346# pfet$140
Xpfet$140_24 vdd vdd m1_5790_24542# m1_3394_25858# pfet$140
Xpfet$140_13 vdd vdd m1_12259_24224# m1_11639_23922# pfet$140
Xpfet$170_1 vdd m1_n4485_20152# vdd m1_n3206_20274# pfet$170
Xpfet$163_0 vdd vdd m1_n7320_25516# m1_n7186_25858# pfet$163
Xnfet$150_4 m1_2912_25858# vss m1_3049_25662# vss nfet$150
Xnfet$153_72 m1_17851_17714# vss m1_18441_17518# vss nfet$153
Xnfet$153_61 m1_20104_16080# vss m1_19747_15778# vss nfet$153
Xnfet$153_50 m1_25747_17714# vss m1_22848_17343# vss nfet$153
Xpfet$142_5 vdd m1_9645_21447# m1_9645_21447# m1_9877_22102# m1_11671_21786# m1_11671_21786#
+ pfet$142
Xpfet$141_104 vdd vdd m1_14127_16080# m1_n7513_20152# pfet$141
Xpfet$146_12 vdd vdd m1_15171_20152# m1_9331_15478# pfet$146
Xpfet$140_2 vdd vdd m1_3394_25858# m1_4509_24346# pfet$140
Xnfet$150_62 m1_24188_23922# vss m1_24808_24224# vss nfet$150
Xnfet$150_51 m1_19644_25858# m1_21729_25658# m1_22522_24542# vss nfet$150
Xnfet$150_40 m1_15598_25662# m1_16442_24224# m1_17546_25658# vss nfet$150
Xnfet$169_27 m1_18310_16080# m1_18310_16080# vss vss m1_19873_17358# vss nfet$169
Xnfet$169_16 m1_19747_15778# m1_19747_15778# m1_19637_18030# m1_19637_18030# m1_19873_17358#
+ vss nfet$169
Xnfet$177_9 m1_n3184_24224# vss m1_n3541_23922# vss nfet$177
Xnfet$150_73 m1_24309_25858# vss m1_21590_21786# vss nfet$150
Xpfet$143_35 vdd m1_n3822_21786# m1_n3822_21786# m1_13373_19850# m1_12935_19550# m1_12935_19550#
+ pfet$143
Xpfet$143_24 vdd m1_n1927_20274# m1_n1927_20274# m1_16890_19850# m1_16452_19550# m1_16452_19550#
+ pfet$143
Xpfet$143_13 vdd m1_n927_19404# m1_n927_19404# m1_n695_19850# m1_n1133_19550# m1_n1133_19550#
+ pfet$143
Xnfet$166_2 m1_31535_19792# m1_32818_20470# vss vss nfet$166
Xnfet$173_3 m1_n6172_16202# m1_n6172_16202# vss vss m1_n6690_16398# vss nfet$173
Xnfet$159_1 m1_n1271_25858# m1_n647_25662# m1_n910_23922# vss nfet$159
Xpfet$158_3 vdd m1_n5461_18030# vdd m1_n6788_16080# pfet$158
Xpfet$165_4 vdd vdd m1_n4485_21904# m1_n3822_21786# pfet$165
Xnfet$152_8 m1_27003_19550# m1_27003_19550# vss vss m1_27441_20470# vss nfet$152
Xpfet$156_0 vdd vdd fout m1_34093_22102# pfet$156
Xpfet$140_69 vdd vdd m1_12875_24346# m1_n7513_20152# pfet$140
Xpfet$140_58 vdd vdd m1_23964_25662# m1_23827_25858# pfet$140
Xpfet$140_47 vdd vdd m1_15943_25858# m1_17058_24346# pfet$140
Xpfet$144_9 vdd vdd m1_22222_21786# m1_21590_21786# pfet$144
Xnfet$171_0 m1_35837_22102# vss m1_n7513_20152# vss nfet$171
Xpfet$140_36 vdd vdd m1_8692_24346# m1_n7513_20152# pfet$140
Xpfet$140_25 vdd vdd m1_4005_21786# m1_3394_25858# pfet$140
Xpfet$140_14 vdd vdd m1_11902_25662# m1_11760_25858# pfet$140
Xpfet$170_2 vdd m1_n5227_20152# vdd m1_n1927_20274# pfet$170
Xpfet$163_1 vdd vdd m1_n6111_25858# m1_n6856_24542# pfet$163
Xnfet$153_73 m1_13668_17714# vss m1_16538_15778# vss nfet$153
Xnfet$153_62 m1_18665_17343# m1_20721_15778# m1_20104_16080# vss nfet$153
Xnfet$153_51 m1_n7513_20152# vss m1_22493_16080# vss nfet$153
Xnfet$150_5 m1_2912_25858# m1_3536_25662# m1_3273_23922# vss nfet$150
Xnfet$153_40 m1_n2250_17343# m1_n194_15778# m1_n811_16080# vss nfet$153
Xpfet$142_6 vdd vdd vdd m1_10505_22402# m1_9288_21786# m1_9288_21786# pfet$142
Xpfet$141_90 vdd m1_19747_15778# m1_18926_16202# m1_18665_17343# pfet$141
Xpfet$146_13 vdd vdd m1_16452_19550# m1_13198_17714# pfet$146
Xpfet$140_3 vdd m1_3394_25858# vdd m1_4997_25658# pfet$140
Xpfet$141_105 vdd vdd m1_14258_17518# m1_13668_17714# pfet$141
Xnfet$169_17 m1_22493_16080# m1_22493_16080# vss vss m1_24056_17358# vss nfet$169
Xnfet$150_74 pd8 vss m1_23356_21786# vss nfet$150
Xnfet$150_63 m1_14556_21786# vss m1_19644_25858# vss nfet$150
Xnfet$150_52 m1_20126_25858# vss m1_22522_24542# vss nfet$150
Xnfet$150_41 pd5 vss m1_12805_21786# vss nfet$150
Xnfet$150_30 m1_n7513_20152# vss m1_17058_24346# vss nfet$150
Xpfet$143_25 vdd vdd vdd m1_17526_19550# m1_13514_15478# m1_13514_15478# pfet$143
Xpfet$143_14 vdd m1_n927_19404# m1_n927_19404# m1_n59_19550# m1_n7383_17599# m1_n7383_17599#
+ pfet$143
Xnfet$166_3 m1_30256_22102# vss m1_32818_21586# vss nfet$166
Xnfet$173_4 m1_28113_15778# m1_28113_15778# m1_28003_18030# m1_28003_18030# m1_28239_17358#
+ vss nfet$173
Xnfet$159_2 m1_n1271_25858# m1_814_25658# m1_1607_24542# vss nfet$159
Xpfet$158_4 vdd vdd m1_26217_17714# m1_26676_16080# pfet$158
Xpfet$165_5 vdd m1_n6839_21786# vdd m1_n5764_21786# pfet$165
Xnfet$152_9 m1_25747_17714# m1_25747_17714# vss vss m1_28073_20470# vss nfet$152
Xnfet$164_0 m1_34843_21786# m1_34843_21786# m1_34093_22102# m1_34093_22102# m1_34329_21430#
+ vss nfet$164
Xpfet$140_59 vdd vdd m1_16322_21786# pd6 pfet$140
Xpfet$140_48 vdd m1_16085_25662# m1_15822_23922# m1_15598_25662# pfet$140
Xpfet$140_37 vdd vdd m1_9973_24542# m1_7577_25858# pfet$140
Xpfet$140_26 vdd m1_4997_25658# m1_5790_24542# m1_3049_25662# pfet$140
Xpfet$140_15 vdd m1_11902_25662# m1_11639_23922# m1_11415_25662# pfet$140
Xpfet$170_3 vdd m1_n6839_20152# vdd m1_n927_19404# pfet$170
Xpfet$149_0 vdd vdd m1_n646_24542# m1_n290_24224# pfet$149
Xnfet$153_74 m1_14482_17343# vss m1_14641_17836# vss nfet$153
Xnfet$153_63 m1_13668_17714# vss m1_14258_17518# vss nfet$153
Xnfet$153_52 m1_23007_17836# m1_24287_16080# m1_23820_18030# vss nfet$153
Xnfet$150_6 m1_3049_25662# m1_3893_24224# m1_4997_25658# vss nfet$150
Xnfet$153_30 sd6 vss m1_5148_15478# vss nfet$153
Xnfet$153_41 m1_n2091_17836# m1_n1168_15778# m1_n1989_16202# vss nfet$153
Xpfet$142_7 vdd m1_354_22513# m1_354_22513# m1_n674_22102# m1_1120_21786# m1_1120_21786#
+ pfet$142
Xpfet$141_91 vdd m1_24287_16080# m1_23820_18030# m1_22848_17343# pfet$141
Xpfet$141_80 vdd vdd m1_15564_15778# m1_15921_16080# pfet$141
Xpfet$146_14 vdd vdd m1_23486_19550# m1_21564_17714# pfet$146
Xpfet$140_4 vdd vdd m1_3893_24224# m1_3273_23922# pfet$140
Xpfet$141_106 vdd vdd m1_14482_17343# m1_17381_17714# pfet$141
Xnfet$169_18 m1_23930_15778# m1_23930_15778# m1_23820_18030# m1_23820_18030# m1_24056_17358#
+ vss nfet$169
Xnfet$150_75 m1_28371_23922# vss m1_28991_24224# vss nfet$150
Xnfet$150_64 m1_19644_25858# vss m1_19781_25662# vss nfet$150
Xnfet$150_53 m1_23827_25858# m1_24451_25662# m1_24188_23922# vss nfet$150
Xnfet$150_42 m1_15943_25858# vss m1_16085_25662# vss nfet$150
Xnfet$150_31 m1_15943_25858# vss m1_18339_24542# vss nfet$150
Xnfet$150_20 pd3 vss m1_5771_21786# vss nfet$150
Xpfet$143_26 vdd m1_n1927_20274# m1_n1927_20274# m1_17526_19550# m1_13198_17714# m1_13198_17714#
+ pfet$143
Xpfet$143_15 vdd vdd vdd m1_n59_19550# m1_n7401_15478# m1_n7401_15478# pfet$143
Xnfet$173_5 m1_26676_16080# m1_26676_16080# vss vss m1_28239_17358# vss nfet$173
Xpfet$158_5 vdd m1_26217_17714# vdd m1_27292_16202# pfet$158
Xnfet$159_3 m1_n1134_25662# m1_n290_24224# m1_814_25658# vss nfet$159
Xpfet$165_6 vdd vdd m1_n6973_21481# m1_n6839_21786# pfet$165
Xnfet$164_1 m1_28490_22513# m1_28490_22513# vss vss m1_34329_21430# vss nfet$164
Xpfet$140_49 vdd m1_20126_25858# vdd m1_21729_25658# pfet$140
Xpfet$140_38 vdd vdd m1_16085_25662# m1_15943_25858# pfet$140
Xpfet$140_27 vdd vdd m1_11278_25858# m1_7522_21786# pfet$140
Xpfet$140_16 vdd vdd m1_5771_21786# pd3 pfet$140
Xnfet$157_0 m1_n3534_17714# vss m1_n6433_17343# vss nfet$157
Xpfet$149_1 vdd m1_n789_25858# vdd m1_814_25658# pfet$149
Xpfet$170_4 vdd vdd m1_n6839_20152# m1_n6973_21481# pfet$170
Xnfet$153_75 sd3 vss m1_17697_15478# vss nfet$153
Xnfet$153_64 m1_13668_17714# vss m1_13198_17714# vss nfet$153
Xnfet$153_53 m1_22848_17343# vss m1_23007_17836# vss nfet$153
Xnfet$150_7 m1_3049_25662# m1_3273_23922# m1_3537_24542# vss nfet$150
Xnfet$153_31 m1_1933_17343# m1_3989_15778# m1_3372_16080# vss nfet$153
Xnfet$153_20 m1_1119_17714# vss m1_1709_17518# vss nfet$153
Xnfet$153_42 m1_n811_16080# vss m1_n1168_15778# vss nfet$153
Xpfet$161_0 vdd vdd vdd m1_n6624_23622# m1_n7082_23622# m1_n7082_23622# pfet$161
Xpfet$142_8 vdd vdd vdd m1_6360_22102# m1_5901_21590# m1_5901_21590# pfet$142
Xpfet$141_92 vdd m1_15454_18030# vdd m1_14127_16080# pfet$141
Xpfet$141_81 vdd vdd m1_13668_17714# m1_14127_16080# pfet$141
Xpfet$141_70 vdd vdd m1_18824_17836# m1_18665_17343# pfet$141
Xpfet$146_15 vdd vdd m1_22205_20152# m1_17697_15478# pfet$146
Xpfet$140_5 vdd m1_3893_24224# m1_4997_25658# m1_2912_25858# pfet$140
Xpfet$141_107 vdd m1_15921_16080# m1_15454_18030# m1_14482_17343# pfet$141
Xnfet$169_19 m1_23109_16202# m1_23109_16202# vss vss m1_22591_16398# vss nfet$169
Xnfet$150_76 m1_28492_25858# vss m1_28634_25662# vss nfet$150
Xnfet$150_65 m1_28492_25858# vss m1_25107_21786# vss nfet$150
Xnfet$150_54 m1_24309_25858# vss m1_24451_25662# vss nfet$150
Xnfet$150_43 m1_15461_25858# vss m1_15598_25662# vss nfet$150
Xnfet$150_32 m1_15461_25858# m1_17546_25658# m1_18339_24542# vss nfet$150
Xnfet$150_21 m1_11278_25858# m1_11902_25662# m1_11639_23922# vss nfet$150
Xnfet$150_10 m1_7577_25858# vss m1_9973_24542# vss nfet$150
Xpfet$143_27 vdd vdd vdd m1_20407_19850# m1_22205_20152# m1_22205_20152# pfet$143
Xpfet$143_16 vdd vdd vdd m1_28077_19550# m1_26063_15478# m1_26063_15478# pfet$143
Xnfet$159_4 m1_32193_25858# m1_34278_25658# m1_35071_24542# vss nfet$159
Xpfet$158_6 vdd vdd m1_28003_18030# m1_28113_15778# pfet$158
Xnfet$173_6 m1_27292_16202# m1_27292_16202# vss vss m1_26774_16398# vss nfet$173
Xpfet$165_7 vdd vdd m1_n6839_21786# m1_n6380_21786# pfet$165
Xnfet$164_2 m1_9645_21447# m1_9645_21447# vss vss m1_30492_21430# vss nfet$164
Xnfet$157_1 m1_n7513_20152# vss m1_n6788_16080# vss nfet$157
Xpfet$140_39 vdd vdd m1_15598_25662# m1_15461_25858# pfet$140
Xpfet$140_28 vdd m1_11639_23922# m1_11903_24542# m1_11278_25858# pfet$140
Xpfet$140_17 vdd vdd m1_7577_25858# m1_8692_24346# pfet$140
Xpfet$149_2 vdd vdd m1_n789_25858# m1_326_24346# pfet$149
Xnfet$150_8 m1_3394_25858# vss m1_3536_25662# vss nfet$150
Xnfet$153_76 m1_14482_17343# m1_16538_15778# m1_15921_16080# vss nfet$153
Xnfet$153_65 m1_14482_17343# m1_14743_16202# m1_14258_17518# vss nfet$153
Xnfet$153_54 m1_22848_17343# m1_23109_16202# m1_22624_17518# vss nfet$153
Xnfet$153_32 m1_2092_17836# m1_3015_15778# m1_2194_16202# vss nfet$153
Xnfet$153_21 m1_1933_17343# m1_2194_16202# m1_1709_17518# vss nfet$153
Xnfet$153_10 m1_11738_16080# vss m1_11381_15778# vss nfet$153
Xnfet$153_43 sd8 vss m1_n3218_15478# vss nfet$153
Xpfet$142_9 vdd m1_3871_22513# m1_3871_22513# m1_3471_22402# m1_4005_21786# m1_4005_21786#
+ pfet$142
Xpfet$154_0 vdd m1_34093_22102# vdd m1_28490_22513# pfet$154
Xpfet$141_93 vdd m1_23820_18030# vdd m1_22493_16080# pfet$141
Xpfet$141_82 vdd m1_13668_17714# vdd m1_14743_16202# pfet$141
Xpfet$141_71 vdd vdd m1_19747_15778# m1_20104_16080# pfet$141
Xpfet$141_60 vdd vdd m1_n194_15778# m1_n3064_17714# pfet$141
Xpfet$161_1 vdd m1_n6856_24542# m1_n6856_24542# m1_n6624_23622# m1_n8283_19850# m1_n8283_19850#
+ pfet$161
Xpfet$141_108 vdd vdd m1_15454_18030# m1_15564_15778# pfet$141
Xpfet$146_16 vdd vdd m1_19969_19550# m1_17381_17714# pfet$146
Xpfet$140_6 vdd vdd m1_3536_25662# m1_3394_25858# pfet$140
Xnfet$150_77 m1_28010_25858# vss m1_28147_25662# vss nfet$150
Xnfet$150_66 m1_28010_25858# m1_30095_25658# m1_30888_24542# vss nfet$150
Xnfet$150_55 m1_23827_25858# vss m1_23964_25662# vss nfet$150
Xnfet$150_44 m1_15822_23922# vss m1_16442_24224# vss nfet$150
Xnfet$150_33 m1_11760_25858# vss m1_14156_24542# vss nfet$150
Xnfet$150_22 m1_11760_25858# vss m1_11902_25662# vss nfet$150
Xnfet$150_11 m1_7522_21786# vss m1_11278_25858# vss nfet$150
Xpfet$143_28 vdd vdd vdd m1_21043_19550# m1_17697_15478# m1_17697_15478# pfet$143
Xpfet$143_17 vdd m1_n3822_20130# m1_n3822_20130# m1_28077_19550# m1_25747_17714# m1_25747_17714#
+ pfet$143
Xnfet$159_5 m1_32330_25662# m1_33174_24224# m1_34278_25658# vss nfet$159
Xnfet$173_7 m1_26676_16080# m1_26676_16080# m1_26217_17714# m1_26217_17714# m1_26774_16398#
+ vss nfet$173
Xpfet$158_7 vdd m1_28003_18030# vdd m1_26676_16080# pfet$158
Xnfet$164_3 m1_7388_22513# m1_7388_22513# m1_30256_22102# m1_30256_22102# m1_30492_21430#
+ vss nfet$164
Xpfet$149_3 vdd m1_n646_24542# vdd m1_326_24346# pfet$149
Xpfet$140_29 vdd vdd m1_11903_24542# m1_12259_24224# pfet$140
Xpfet$140_18 vdd vdd m1_11415_25662# m1_11278_25858# pfet$140
Xnfet$157_2 m1_n4994_16080# vss m1_n5351_15778# vss nfet$157
Xnfet$150_9 m1_3273_23922# vss m1_3893_24224# vss nfet$150
Xnfet$153_77 sd4 vss m1_13514_15478# vss nfet$153
Xnfet$153_66 m1_n7513_20152# vss m1_14127_16080# vss nfet$153
Xnfet$153_55 m1_22034_17714# vss m1_24904_15778# vss nfet$153
Xnfet$153_44 m1_n2091_17836# m1_n811_16080# m1_n1278_18030# vss nfet$153
Xnfet$153_33 sd7 vss m1_965_15478# vss nfet$153
Xnfet$153_22 m1_6116_17343# m1_6377_16202# m1_5892_17518# vss nfet$153
Xnfet$153_11 m1_10299_17343# m1_12355_15778# m1_11738_16080# vss nfet$153
Xnfet$162_0 m1_11039_21786# m1_11039_21786# vss vss m1_9877_21586# vss nfet$162
Xpfet$154_1 vdd vdd m1_34093_22102# m1_34843_21786# pfet$154
Xpfet$141_94 vdd vdd m1_22624_17518# m1_22034_17714# pfet$141
Xpfet$141_83 vdd m1_16538_15778# m1_15921_16080# m1_14641_17836# pfet$141
Xpfet$141_72 vdd m1_20721_15778# m1_20104_16080# m1_18824_17836# pfet$141
Xpfet$141_61 vdd m1_n811_16080# m1_n1278_18030# m1_n2250_17343# pfet$141
Xpfet$141_50 vdd m1_n1168_15778# m1_n1989_16202# m1_n2250_17343# pfet$141
Xpfet$147_0 vdd vdd m1_n7401_15478# sd9 pfet$147
Xpfet$141_109 vdd vdd m1_10299_17343# m1_13198_17714# pfet$141
Xpfet$146_17 vdd vdd m1_25722_20152# m1_21880_15478# pfet$146
Xpfet$140_7 vdd vdd m1_7232_25662# m1_7095_25858# pfet$140
Xnfet$150_78 m1_28010_25858# m1_28634_25662# m1_28371_23922# vss nfet$150
Xnfet$150_67 m1_28492_25858# vss m1_30888_24542# vss nfet$150
Xnfet$150_56 m1_19781_25662# m1_20625_24224# m1_21729_25658# vss nfet$150
Xnfet$150_45 m1_15461_25858# m1_16085_25662# m1_15822_23922# vss nfet$150
Xnfet$150_34 m1_11278_25858# m1_13363_25658# m1_14156_24542# vss nfet$150
Xnfet$150_23 m1_11278_25858# vss m1_11415_25662# vss nfet$150
Xnfet$150_12 m1_7577_25858# vss m1_7522_21786# vss nfet$150
Xpfet$143_29 vdd vdd vdd m1_23924_19850# m1_25722_20152# m1_25722_20152# pfet$143
Xpfet$143_18 vdd vdd vdd m1_27441_19850# m1_29239_20152# m1_29239_20152# pfet$143
Xnfet$159_6 m1_32193_25858# m1_32817_25662# m1_32554_23922# vss nfet$159
Xpfet$149_4 vdd vdd m1_32675_25947# m1_33790_24346# pfet$149
Xpfet$140_19 vdd vdd m1_7095_25858# m1_4005_21786# pfet$140
Xnfet$157_3 m1_n6433_17343# vss m1_n6274_17836# vss nfet$157
Xnfet$153_78 m1_14641_17836# m1_15564_15778# m1_14743_16202# vss nfet$153
Xnfet$153_67 m1_17381_17714# vss m1_14482_17343# vss nfet$153
Xnfet$153_56 m1_24287_16080# vss m1_23930_15778# vss nfet$153
Xnfet$153_45 m1_n3064_17714# vss m1_n194_15778# vss nfet$153
Xnfet$155_0 m1_n3534_17714# vss m1_2384_19550# vss nfet$155
Xnfet$153_34 m1_n2250_17343# vss m1_n2091_17836# vss nfet$153
Xnfet$153_23 m1_5302_17714# vss m1_4832_17714# vss nfet$153
Xnfet$153_12 m1_9485_17714# vss m1_12355_15778# vss nfet$153
Xnfet$162_1 m1_11671_21786# m1_11671_21786# vss vss m1_10509_21586# vss nfet$162
Xpfet$154_2 vdd vdd m1_30256_22102# m1_7388_22513# pfet$154
Xpfet$147_1 vdd vdd m1_21880_15478# sd2 pfet$147
Xpfet$141_95 vdd vdd m1_21564_17714# m1_22034_17714# pfet$141
Xpfet$141_84 vdd vdd m1_17381_17714# m1_17851_17714# pfet$141
Xpfet$141_73 vdd vdd m1_16538_15778# m1_13668_17714# pfet$141
Xpfet$141_62 vdd vdd m1_23007_17836# m1_22848_17343# pfet$141
Xpfet$141_40 vdd m1_10560_16202# m1_10075_17518# m1_10458_17836# pfet$141
Xpfet$141_51 vdd vdd m1_n1168_15778# m1_n811_16080# pfet$141
Xpfet$140_8 vdd vdd m1_8076_24224# m1_7456_23922# pfet$140
Xpfet$140_110 vdd m1_11903_24542# vdd m1_12875_24346# pfet$140
Xnfet$150_79 pd7 vss m1_19839_21786# vss nfet$150
Xnfet$150_68 m1_n7513_20152# vss m1_29607_24346# vss nfet$150
Xnfet$150_57 m1_20126_25858# vss m1_20268_25662# vss nfet$150
Xnfet$150_46 m1_20126_25858# vss m1_18073_21786# vss nfet$150
Xnfet$150_35 m1_15598_25662# m1_15822_23922# m1_16086_24542# vss nfet$150
Xnfet$150_24 m1_7095_25858# m1_7719_25662# m1_7456_23922# vss nfet$150
Xnfet$150_13 m1_11415_25662# m1_11639_23922# m1_11903_24542# vss nfet$150
Xpfet$143_19 vdd m1_n3822_20130# m1_n3822_20130# m1_27441_19850# m1_27003_19550# m1_27003_19550#
+ pfet$143
Xnfet$159_7 m1_32330_25662# m1_32554_23922# m1_32818_24542# vss nfet$159
Xnfet$185_0 m1_n6839_20152# vss m1_n8145_21908# vss nfet$185
Xnfet$157_4 m1_n7247_17714# vss m1_n4377_15778# vss nfet$157
Xpfet$149_5 vdd m1_32675_25947# vdd m1_34278_25658# pfet$149
Xnfet$153_79 m1_15921_16080# vss m1_15564_15778# vss nfet$153
Xnfet$153_68 m1_18665_17343# m1_18926_16202# m1_18441_17518# vss nfet$153
Xnfet$153_57 m1_22848_17343# m1_24904_15778# m1_24287_16080# vss nfet$153
Xnfet$153_46 m1_22034_17714# vss m1_21564_17714# vss nfet$153
Xnfet$153_24 m1_4832_17714# vss m1_1933_17343# vss nfet$153
Xnfet$153_13 m1_10458_17836# m1_11381_15778# m1_10560_16202# vss nfet$153
Xnfet$153_35 m1_n7513_20152# vss m1_5761_16080# vss nfet$153
Xpfet$147_2 vdd vdd m1_26063_15478# sd1 pfet$147
Xpfet$154_3 vdd m1_31535_22102# vdd m1_3871_22513# pfet$154
Xnfet$155_1 m1_n3218_15478# vss m1_4620_20152# vss nfet$155
Xnfet$162_2 m1_8154_21786# m1_8154_21786# vss vss m1_6992_21586# vss nfet$162
Xpfet$141_96 vdd vdd m1_18665_17343# m1_21564_17714# pfet$141
Xpfet$141_85 vdd m1_18926_16202# m1_18441_17518# m1_18824_17836# pfet$141
Xpfet$141_74 vdd vdd m1_14641_17836# m1_14482_17343# pfet$141
Xpfet$141_63 vdd m1_23930_15778# m1_23109_16202# m1_22848_17343# pfet$141
Xpfet$141_30 vdd vdd m1_1933_17343# m1_4832_17714# pfet$141
Xpfet$141_41 vdd vdd m1_10075_17518# m1_9485_17714# pfet$141
Xpfet$141_52 vdd m1_n3064_17714# vdd m1_n1989_16202# pfet$141
Xpfet$140_9 vdd m1_7719_25662# m1_7456_23922# m1_7232_25662# pfet$140
Xpfet$152_0 vdd m1_n647_25662# m1_n910_23922# m1_n1134_25662# pfet$152
Xpfet$140_100 vdd vdd m1_29607_24346# m1_n7513_20152# pfet$140
Xnfet$150_69 m1_24309_25858# vss m1_26705_24542# vss nfet$150
Xnfet$150_58 m1_20005_23922# vss m1_20625_24224# vss nfet$150
Xnfet$150_47 m1_23964_25662# m1_24188_23922# m1_24452_24542# vss nfet$150
Xnfet$150_36 m1_11760_25858# vss m1_11039_21786# vss nfet$150
Xnfet$150_25 m1_7232_25662# m1_8076_24224# m1_9180_25658# vss nfet$150
Xnfet$150_14 m1_n7513_20152# vss m1_8692_24346# vss nfet$150
Xnfet$178_0 m1_n9952_24224# m1_n9952_24224# m1_n10308_24542# m1_n10308_24542# m1_n9854_24542#
+ vss nfet$178
Xnfet$157_5 m1_n7247_17714# vss m1_n6657_17518# vss nfet$157
Xpfet$149_6 vdd vdd m1_32818_24542# m1_33174_24224# pfet$149
Xnfet$153_69 m1_17851_17714# vss m1_17381_17714# vss nfet$153
Xnfet$153_58 m1_23007_17836# m1_23930_15778# m1_23109_16202# vss nfet$153
Xnfet$153_47 m1_22034_17714# vss m1_22624_17518# vss nfet$153
Xnfet$153_25 m1_2092_17836# m1_3372_16080# m1_2905_18030# vss nfet$153
Xnfet$153_14 m1_6116_17343# m1_8172_15778# m1_7555_16080# vss nfet$153
Xnfet$153_36 m1_n3064_17714# vss m1_n2474_17518# vss nfet$153
Xpfet$154_4 vdd m1_30256_22102# vdd m1_9645_21447# pfet$154
Xnfet$155_2 m1_n7401_15478# vss m1_1103_20152# vss nfet$155
Xnfet$162_3 m1_7522_21786# m1_7522_21786# vss vss m1_6360_21586# vss nfet$162
Xpfet$141_97 vdd vdd m1_22493_16080# m1_n7513_20152# pfet$141
Xpfet$141_86 vdd m1_19637_18030# vdd m1_18310_16080# pfet$141
Xpfet$141_75 vdd vdd m1_17697_15478# sd3 pfet$141
Xpfet$141_64 vdd vdd m1_23930_15778# m1_24287_16080# pfet$141
Xpfet$141_20 vdd vdd m1_1119_17714# m1_1578_16080# pfet$141
Xpfet$141_31 vdd m1_3372_16080# m1_2905_18030# m1_1933_17343# pfet$141
Xpfet$141_42 vdd m1_11271_18030# vdd m1_9944_16080# pfet$141
Xpfet$141_53 vdd vdd m1_n3218_15478# sd8 pfet$141
Xnfet$160_0 pd1 vss m1_n1263_21786# vss nfet$160
Xpfet$145_0 vdd vdd m1_n6274_17836# m1_n6433_17343# pfet$145
Xpfet$152_1 vdd m1_n910_23922# m1_n646_24542# m1_n1271_25858# pfet$152
Xpfet$140_101 vdd vdd m1_28010_25858# m1_21590_21786# pfet$140
Xnfet$150_59 m1_19644_25858# m1_20268_25662# m1_20005_23922# vss nfet$150
Xnfet$150_48 m1_18073_21786# vss m1_23827_25858# vss nfet$150
Xnfet$150_37 m1_11039_21786# vss m1_15461_25858# vss nfet$150
Xnfet$150_26 m1_7095_25858# m1_9180_25658# m1_9973_24542# vss nfet$150
Xnfet$150_15 m1_7232_25662# m1_7456_23922# m1_7720_24542# vss nfet$150
Xnfet$178_1 m1_n9336_24346# m1_n9336_24346# m1_n8625_26174# m1_n8625_26174# m1_n8389_25502#
+ vss nfet$178
Xnfet$157_6 m1_n7247_17714# vss m1_n7383_17599# vss nfet$157
Xpfet$149_7 vdd m1_32818_24542# vdd m1_33790_24346# pfet$149
Xnfet$153_59 m1_17851_17714# vss m1_20721_15778# vss nfet$153
Xnfet$153_48 m1_18824_17836# m1_20104_16080# m1_19637_18030# vss nfet$153
Xnfet$155_3 m1_649_17714# vss m1_5901_19550# vss nfet$155
Xnfet$153_26 m1_5302_17714# vss m1_5892_17518# vss nfet$153
Xnfet$153_15 m1_5302_17714# vss m1_8172_15778# vss nfet$153
Xnfet$153_37 m1_n7513_20152# vss m1_n2605_16080# vss nfet$153
Xnfet$162_4 m1_1120_21786# m1_1120_21786# vss vss m1_n42_21586# vss nfet$162
Xpfet$141_98 vdd m1_20104_16080# m1_19637_18030# m1_18665_17343# pfet$141
Xpfet$141_87 vdd vdd m1_18310_16080# m1_n7513_20152# pfet$141
Xpfet$141_76 vdd m1_17851_17714# vdd m1_18926_16202# pfet$141
Xpfet$141_65 vdd m1_24904_15778# m1_24287_16080# m1_23007_17836# pfet$141
Xpfet$141_21 vdd vdd m1_965_15478# sd7 pfet$141
Xpfet$141_10 vdd m1_8172_15778# m1_7555_16080# m1_6275_17836# pfet$141
Xpfet$141_32 vdd vdd m1_2905_18030# m1_3015_15778# pfet$141
Xpfet$141_43 vdd vdd m1_11271_18030# m1_11381_15778# pfet$141
Xpfet$141_54 vdd vdd m1_n1278_18030# m1_n1168_15778# pfet$141
Xnfet$160_1 pd2 vss m1_2254_21786# vss nfet$160
Xnfet$153_0 m1_9485_17714# vss m1_9015_17714# vss nfet$153
Xpfet$145_1 vdd vdd m1_n4377_15778# m1_n7247_17714# pfet$145
Xpfet$152_2 vdd m1_n290_24224# m1_814_25658# m1_n1271_25858# pfet$152
Xpfet$140_102 vdd m1_28371_23922# m1_28635_24542# m1_28010_25858# pfet$140
Xnfet$150_49 m1_19781_25662# m1_20005_23922# m1_20269_24542# vss nfet$150
Xnfet$150_38 m1_n7513_20152# vss m1_12875_24346# vss nfet$150
Xnfet$150_27 m1_7577_25858# vss m1_7719_25662# vss nfet$150
Xnfet$150_16 m1_4005_21786# vss m1_7095_25858# vss nfet$150
Xnfet$178_2 m1_n8848_25658# m1_n8848_25658# vss vss m1_n8389_25502# vss nfet$178
Xpfet$144_10 vdd vdd m1_23486_21590# m1_23356_21786# pfet$144
Xnfet$157_7 m1_26217_17714# vss m1_26807_17518# vss nfet$157
Xnfet$183_0 m1_n927_19404# m1_n927_19404# vss vss m1_n6282_20470# vss nfet$183
Xpfet$168_0 vdd vdd vdd m1_n8047_19550# m1_n7513_20152# m1_n7513_20152# pfet$168
Xnfet$153_49 m1_21564_17714# vss m1_18665_17343# vss nfet$153
Xnfet$155_4 m1_4832_17714# vss m1_9418_19550# vss nfet$155
Xnfet$153_27 m1_1119_17714# vss m1_3989_15778# vss nfet$153
Xnfet$153_16 m1_6275_17836# m1_7198_15778# m1_6377_16202# vss nfet$153
Xnfet$153_38 m1_n2250_17343# m1_n1989_16202# m1_n2474_17518# vss nfet$153
Xnfet$162_5 m1_4005_21786# m1_4005_21786# vss vss m1_2843_21586# vss nfet$162
Xpfet$141_99 vdd m1_23109_16202# m1_22624_17518# m1_23007_17836# pfet$141
Xpfet$141_88 vdd vdd m1_18441_17518# m1_17851_17714# pfet$141
Xpfet$141_77 vdd vdd m1_17851_17714# m1_18310_16080# pfet$141
Xpfet$141_66 vdd vdd m1_24904_15778# m1_22034_17714# pfet$141
Xpfet$141_22 vdd vdd m1_3015_15778# m1_3372_16080# pfet$141
Xpfet$141_11 vdd vdd m1_9485_17714# m1_9944_16080# pfet$141
Xpfet$141_33 vdd vdd m1_5892_17518# m1_5302_17714# pfet$141
Xpfet$141_44 vdd vdd m1_649_17714# m1_1119_17714# pfet$141
Xpfet$141_55 vdd vdd m1_n2474_17518# m1_n3064_17714# pfet$141
Xnfet$160_2 pd9 vss m1_26873_21786# vss nfet$160
Xnfet$153_1 m1_9015_17714# vss m1_6116_17343# vss nfet$153
Xpfet$140_103 vdd vdd m1_28635_24542# m1_28991_24224# pfet$140
Xnfet$150_39 pd4 vss m1_9288_21786# vss nfet$150
Xpfet$152_3 vdd m1_814_25658# m1_1607_24542# m1_n1134_25662# pfet$152
Xnfet$150_28 m1_3394_25858# vss m1_4005_21786# vss nfet$150
Xnfet$150_17 m1_11639_23922# vss m1_12259_24224# vss nfet$150
Xpfet$145_2 vdd vdd m1_n5351_15778# m1_n4994_16080# pfet$145
Xpfet$150_0 vdd vdd vdd m1_33050_22344# m1_31535_22102# m1_31535_22102# pfet$150
Xnfet$178_3 m1_n9336_24346# m1_n9336_24346# vss vss m1_n9854_24542# vss nfet$178
Xpfet$144_11 vdd vdd m1_18705_21786# m1_18073_21786# pfet$144
Xnfet$157_8 m1_n7513_20152# vss m1_26676_16080# vss nfet$157
Xnfet$176_0 m1_n3822_20130# m1_n3822_20130# m1_n4485_20152# m1_n4485_20152# m1_n3724_20470#
+ vss nfet$176
Xnfet$183_1 m1_n2543_20130# m1_n2543_20130# m1_n5227_20152# m1_n5227_20152# m1_n2445_20470#
+ vss nfet$183
Xpfet$168_1 vdd m1_n8283_19850# m1_n8283_19850# m1_n8047_19550# m1_n8283_20611# m1_n8283_20611#
+ pfet$168
Xnfet$155_5 m1_965_15478# vss m1_8137_20152# vss nfet$155
Xnfet$153_28 m1_1933_17343# vss m1_2092_17836# vss nfet$153
Xnfet$153_17 m1_649_17714# vss m1_n2250_17343# vss nfet$153
Xnfet$153_39 m1_n3064_17714# vss m1_n3534_17714# vss nfet$153
Xnfet$162_6 m1_4637_21786# m1_4637_21786# vss vss m1_3475_21586# vss nfet$162
Xpfet$141_12 vdd m1_3989_15778# m1_3372_16080# m1_2092_17836# pfet$141
Xpfet$141_89 vdd vdd m1_22848_17343# m1_25747_17714# pfet$141
Xpfet$141_78 vdd vdd m1_13514_15478# sd4 pfet$141
Xpfet$141_67 vdd m1_22034_17714# vdd m1_23109_16202# pfet$141
Xpfet$141_23 vdd m1_5302_17714# vdd m1_6377_16202# pfet$141
Xpfet$141_34 vdd vdd m1_5761_16080# m1_n7513_20152# pfet$141
Xpfet$141_45 vdd vdd m1_9944_16080# m1_n7513_20152# pfet$141
Xpfet$141_56 vdd m1_n1278_18030# vdd m1_n2605_16080# pfet$141
Xnfet$153_2 m1_6275_17836# m1_7555_16080# m1_7088_18030# vss nfet$153
Xpfet$152_4 vdd m1_33174_24224# m1_34278_25658# m1_32193_25858# pfet$152
Xpfet$145_3 vdd vdd m1_n6657_17518# m1_n7247_17714# pfet$145
Xpfet$140_104 vdd m1_25912_25658# m1_26705_24542# m1_23964_25662# pfet$140
Xnfet$150_29 m1_15943_25858# vss m1_14556_21786# vss nfet$150
Xnfet$150_18 m1_7095_25858# vss m1_7232_25662# vss nfet$150
Xpfet$143_0 vdd m1_2590_19404# m1_2590_19404# m1_3458_19550# m1_n3534_17714# m1_n3534_17714#
+ pfet$143
Xnfet$178_4 m1_n4978_24224# m1_n4978_24224# m1_n10452_25858# m1_n10452_25858# m1_n4880_24542#
+ vss nfet$178
Xpfet$144_12 vdd vdd m1_16452_21590# m1_16322_21786# pfet$144
Xnfet$157_9 m1_n10452_25858# vss m1_27031_17343# vss nfet$157
Xnfet$169_0 m1_7198_15778# m1_7198_15778# m1_7088_18030# m1_7088_18030# m1_7324_17358#
+ vss nfet$169
Xnfet$176_1 m1_n1927_20274# m1_n1927_20274# vss vss m1_n2445_20470# vss nfet$176
Xpfet$168_2 vdd m1_n8283_20611# m1_n8283_20611# m1_n8047_22344# m1_n8145_21908# m1_n8145_21908#
+ pfet$168
Xnfet$153_29 m1_3372_16080# vss m1_3015_15778# vss nfet$153
Xnfet$153_18 m1_1119_17714# vss m1_649_17714# vss nfet$153
Xnfet$162_7 m1_488_21786# m1_488_21786# vss vss m1_n674_21586# vss nfet$162
Xnfet$155_6 m1_9015_17714# vss m1_12935_19550# vss nfet$155
Xpfet$141_79 vdd m1_15564_15778# m1_14743_16202# m1_14482_17343# pfet$141
Xpfet$141_68 vdd vdd m1_22034_17714# m1_22493_16080# pfet$141
Xpfet$141_13 vdd vdd m1_5148_15478# sd6 pfet$141
Xpfet$141_24 vdd m1_6377_16202# m1_5892_17518# m1_6275_17836# pfet$141
Xpfet$141_35 vdd vdd m1_9015_17714# m1_9485_17714# pfet$141
Xpfet$141_46 vdd vdd m1_n2250_17343# m1_649_17714# pfet$141
Xpfet$141_57 vdd m1_n1989_16202# m1_n2474_17518# m1_n2091_17836# pfet$141
Xpfet$166_10 vdd vdd m1_n10933_25858# fin pfet$166
Xnfet$153_3 m1_n7513_20152# vss m1_9944_16080# vss nfet$153
Xpfet$152_5 vdd m1_32817_25662# m1_32554_23922# m1_32330_25662# pfet$152
Xpfet$145_4 vdd vdd m1_n6433_17343# m1_n3534_17714# pfet$145
Xpfet$140_105 vdd vdd m1_30888_24542# m1_28492_25858# pfet$140
Xnfet$150_19 m1_7456_23922# vss m1_8076_24224# vss nfet$150
Xnfet$151_0 m1_n1133_21590# m1_n1133_21590# m1_354_22513# m1_354_22513# m1_n674_21586#
+ vss nfet$151
Xpfet$143_1 vdd vdd vdd m1_2822_19850# m1_4620_20152# m1_4620_20152# pfet$143
Xnfet$178_5 m1_n4362_24346# m1_n4362_24346# vss vss m1_n4880_24542# vss nfet$178
Xpfet$144_13 vdd vdd m1_15188_21786# m1_14556_21786# pfet$144
Xnfet$169_1 m1_5761_16080# m1_5761_16080# vss vss m1_7324_17358# vss nfet$169
Xnfet$176_2 m1_n3206_20274# m1_n3206_20274# vss vss m1_n3724_20470# vss nfet$176
Xnfet$153_19 m1_n7513_20152# vss m1_1578_16080# vss nfet$153
Xpfet$168_3 vdd vdd vdd m1_n8047_22344# m1_n8283_19850# m1_n8283_19850# pfet$168
Xnfet$162_8 m1_25739_21786# m1_25739_21786# vss vss m1_24577_21586# vss nfet$162
Xnfet$155_7 m1_5148_15478# vss m1_11654_20152# vss nfet$155
Xnfet$181_0 m1_n8283_20611# vss m1_n8283_19850# vss nfet$181
Xpfet$141_69 vdd vdd m1_20721_15778# m1_17851_17714# pfet$141
Xpfet$141_14 vdd vdd m1_2092_17836# m1_1933_17343# pfet$141
Xpfet$141_25 vdd vdd m1_1709_17518# m1_1119_17714# pfet$141
Xpfet$141_36 vdd vdd m1_6116_17343# m1_9015_17714# pfet$141
Xpfet$141_47 vdd m1_11738_16080# m1_11271_18030# m1_10299_17343# pfet$141
Xpfet$141_58 vdd vdd m1_n3534_17714# m1_n3064_17714# pfet$141
Xpfet$166_0 vdd vdd m1_n10796_25662# m1_n10933_25858# pfet$166
Xpfet$166_11 vdd vdd m1_n9336_24346# vss pfet$166
Xnfet$153_4 m1_10299_17343# m1_10560_16202# m1_10075_17518# vss nfet$153
Xpfet$152_6 vdd m1_34278_25658# m1_35071_24542# m1_32330_25662# pfet$152
Xpfet$145_5 vdd vdd m1_n6788_16080# m1_n7513_20152# pfet$145
Xpfet$140_106 vdd vdd m1_25107_21786# m1_28492_25858# pfet$140
Xnfet$151_1 m1_n1263_21786# m1_n1263_21786# m1_354_22513# m1_354_22513# m1_n42_21586#
+ vss nfet$151
Xpfet$143_2 vdd m1_2590_19404# m1_2590_19404# m1_2822_19850# m1_2384_19550# m1_2384_19550#
+ pfet$143
Xnfet$178_6 m1_n4978_24224# m1_n4978_24224# vss vss m1_n3415_25502# vss nfet$178
Xpfet$144_14 vdd vdd m1_19969_21590# m1_19839_21786# pfet$144
Xnfet$169_2 m1_9944_16080# m1_9944_16080# vss vss m1_11507_17358# vss nfet$169
Xnfet$176_3 m1_n6973_21481# m1_n6973_21481# m1_n6839_20152# m1_n6839_20152# m1_n6282_20470#
+ vss nfet$176
Xnfet$162_9 m1_25107_21786# m1_25107_21786# vss vss m1_23945_21586# vss nfet$162
Xnfet$155_8 m1_n7383_17599# vss m1_n1133_19550# vss nfet$155
Xpfet$141_15 vdd vdd m1_5302_17714# m1_5761_16080# pfet$141
Xpfet$141_26 vdd vdd m1_4832_17714# m1_5302_17714# pfet$141
Xpfet$141_37 vdd m1_7555_16080# m1_7088_18030# m1_6116_17343# pfet$141
Xpfet$141_48 vdd vdd m1_n3064_17714# m1_n2605_16080# pfet$141
Xnfet$181_1 m1_n7513_20152# m1_n8283_19850# vss vss nfet$181
Xpfet$141_59 vdd vdd m1_n2605_16080# m1_n7513_20152# pfet$141
Xpfet$166_1 vdd vdd m1_n10309_25662# m1_n10452_25858# pfet$166
Xnfet$174_0 m1_n10452_25858# m1_n10452_25858# m1_n7186_25858# m1_n7186_25858# m1_n6629_25502#
+ vss nfet$174
Xpfet$159_0 vdd m1_n4377_15778# m1_n4994_16080# m1_n6274_17836# pfet$159
Xpfet$166_12 vdd vdd m1_n7082_23622# m1_n8625_26174# pfet$166
Xpfet$152_7 vdd m1_32554_23922# m1_32818_24542# m1_32193_25858# pfet$152
Xnfet$153_5 m1_10458_17836# m1_11738_16080# m1_11271_18030# vss nfet$153
Xpfet$145_6 vdd vdd m1_n7383_17599# m1_n7247_17714# pfet$145
Xpfet$140_107 vdd m1_24309_25858# vdd m1_25912_25658# pfet$140
Xnfet$151_2 m1_9288_21786# m1_9288_21786# m1_9645_21447# m1_9645_21447# m1_10509_21586#
+ vss nfet$151
Xpfet$143_3 vdd vdd vdd m1_3458_19550# m1_n3218_15478# m1_n3218_15478# pfet$143
Xpfet$141_0 vdd vdd m1_12355_15778# m1_9485_17714# pfet$141
Xnfet$178_7 m1_n3541_23922# m1_n3541_23922# m1_n3651_26174# m1_n3651_26174# m1_n3415_25502#
+ vss nfet$178
Xpfet$144_15 vdd vdd m1_27003_21590# m1_26873_21786# pfet$144
Xnfet$169_3 m1_11381_15778# m1_11381_15778# m1_11271_18030# m1_11271_18030# m1_11507_17358#
+ vss nfet$169
Xnfet$176_4 m1_2590_19404# m1_2590_19404# vss vss m1_n2445_21430# vss nfet$176
Xnfet$155_9 m1_25747_17714# vss m1_27003_19550# vss nfet$155
Xnfet$167_0 m1_34093_22102# vss fout vss nfet$167
Xpfet$141_16 vdd vdd m1_3989_15778# m1_1119_17714# pfet$141
Xpfet$141_27 vdd m1_2194_16202# m1_1709_17518# m1_2092_17836# pfet$141
Xpfet$141_38 vdd vdd m1_7088_18030# m1_7198_15778# pfet$141
Xpfet$141_49 vdd m1_n194_15778# m1_n811_16080# m1_n2091_17836# pfet$141
Xnfet$181_2 m1_n8145_21908# vss m1_n8283_20611# vss nfet$181
Xnfet$174_1 m1_n6111_25858# m1_n6111_25858# vss vss m1_n6629_25502# vss nfet$174
Xpfet$159_1 vdd m1_n5351_15778# m1_n6172_16202# m1_n6433_17343# pfet$159
Xpfet$166_2 vdd vdd m1_n9952_24224# m1_n10572_23922# pfet$166
Xpfet$166_13 vdd vdd m1_n8055_24542# m1_n8625_26174# pfet$166
Xnfet$153_6 m1_6116_17343# vss m1_6275_17836# vss nfet$153
Xpfet$140_108 vdd vdd m1_25424_24346# m1_n7513_20152# pfet$140
Xpfet$145_7 vdd vdd m1_27190_17836# m1_27031_17343# pfet$145
Xpfet$171_0 vdd vdd vdd m1_n5019_19550# m1_n4485_20152# m1_n4485_20152# pfet$171
Xnfet$149_20 m1_21241_24346# m1_21241_24346# m1_20126_25858# m1_20126_25858# m1_22188_25502#
+ vss nfet$149
Xpfet$143_4 vdd m1_6107_19404# m1_6107_19404# m1_6339_19850# m1_5901_19550# m1_5901_19550#
+ pfet$143
Xnfet$151_3 m1_9418_21590# m1_9418_21590# m1_9645_21447# m1_9645_21447# m1_9877_21586#
+ vss nfet$151
Xnfet$151_10 m1_19839_21786# m1_19839_21786# m1_21456_22513# m1_21456_22513# m1_21060_21586#
+ vss nfet$151
Xpfet$141_1 vdd vdd m1_11381_15778# m1_11738_16080# pfet$141
Xpfet$144_16 vdd vdd m1_29256_21786# m1_28624_21786# pfet$144
Xnfet$176_5 m1_6107_19404# m1_6107_19404# m1_n5227_21418# m1_n5227_21418# m1_n2445_21430#
+ vss nfet$176
Xnfet$169_4 m1_10560_16202# m1_10560_16202# vss vss m1_10042_16398# vss nfet$169
Xpfet$141_17 vdd vdd m1_n2091_17836# m1_n2250_17343# pfet$141
Xnfet$181_3 m1_n8283_19850# m1_n8283_20611# vss vss nfet$181
Xpfet$141_28 vdd m1_2905_18030# vdd m1_1578_16080# pfet$141
Xpfet$141_39 vdd m1_7088_18030# vdd m1_5761_16080# pfet$141
Xpfet$159_2 vdd m1_n4994_16080# m1_n5461_18030# m1_n6433_17343# pfet$159
Xpfet$166_3 vdd vdd m1_n4978_24224# vss pfet$166
Xnfet$154_10 m1_21590_21786# vss m1_22222_21786# vss nfet$154
Xnfet$153_7 m1_9485_17714# vss m1_10075_17518# vss nfet$153
Xpfet$145_8 vdd vdd m1_28113_15778# m1_28470_16080# pfet$145
Xpfet$140_109 vdd m1_12259_24224# m1_13363_25658# m1_11278_25858# pfet$140
Xpfet$164_0 vdd vdd m1_n8625_26174# m1_n9336_24346# pfet$164
Xnfet$149_21 m1_28991_24224# m1_28991_24224# m1_28635_24542# m1_28635_24542# m1_29089_24542#
+ vss nfet$149
Xnfet$149_10 m1_17546_25658# m1_17546_25658# vss vss m1_18005_25502# vss nfet$149
Xpfet$143_5 vdd vdd vdd m1_n695_19850# m1_1103_20152# m1_1103_20152# pfet$143
Xnfet$151_4 m1_5901_21590# m1_5901_21590# m1_7388_22513# m1_7388_22513# m1_6360_21586#
+ vss nfet$151
Xnfet$151_11 m1_19969_21590# m1_19969_21590# m1_21456_22513# m1_21456_22513# m1_20428_21586#
+ vss nfet$151
Xpfet$141_2 vdd m1_12355_15778# m1_11738_16080# m1_10458_17836# pfet$141
Xpfet$144_17 vdd vdd m1_25739_21786# m1_25107_21786# pfet$144
Xnfet$162_10 m1_21590_21786# m1_21590_21786# vss vss m1_20428_21586# vss nfet$162
Xnfet$157_10 m1_26217_17714# vss m1_29087_15778# vss nfet$157
Xnfet$169_5 m1_9944_16080# m1_9944_16080# m1_9485_17714# m1_9485_17714# m1_10042_16398#
+ vss nfet$169
Xnfet$176_6 m1_n5764_21786# m1_n5764_21786# vss vss m1_n6282_21430# vss nfet$176
Xpfet$141_18 vdd m1_1119_17714# vdd m1_2194_16202# pfet$141
Xpfet$141_29 vdd vdd m1_1578_16080# m1_n7513_20152# pfet$141
Xpfet$159_3 vdd m1_n6172_16202# m1_n6657_17518# m1_n6274_17836# pfet$159
Xpfet$166_4 vdd vdd m1_n5571_25662# m1_n10452_25858# pfet$166
Xnfet$153_8 m1_7555_16080# vss m1_7198_15778# vss nfet$153
Xnfet$154_11 m1_18073_21786# vss m1_18705_21786# vss nfet$154
Xnfet$170_10 m1_9331_15478# m1_9331_15478# m1_n3822_21786# m1_n3822_21786# m1_13373_20470#
+ vss nfet$170
Xpfet$145_9 vdd vdd m1_29087_15778# m1_26217_17714# pfet$145
Xnfet$172_0 m1_n6274_17836# m1_n4994_16080# m1_n5461_18030# vss nfet$172
Xpfet$157_0 vdd m1_32818_20470# m1_32818_20470# m1_33050_19550# m1_30256_19792# m1_30256_19792#
+ pfet$157
Xpfet$164_1 vdd m1_n8625_26174# vdd m1_n8848_25658# pfet$164
Xnfet$149_22 m1_29607_24346# m1_29607_24346# vss vss m1_29089_24542# vss nfet$149
Xnfet$149_11 m1_16442_24224# m1_16442_24224# m1_16086_24542# m1_16086_24542# m1_16540_24542#
+ vss nfet$149
Xnfet$151_5 m1_2254_21786# m1_2254_21786# m1_3871_22513# m1_3871_22513# m1_3475_21586#
+ vss nfet$151
Xpfet$143_6 vdd vdd vdd m1_6339_19850# m1_8137_20152# m1_8137_20152# pfet$143
Xnfet$151_12 m1_16322_21786# m1_16322_21786# m1_17939_22513# m1_17939_22513# m1_17543_21586#
+ vss nfet$151
Xpfet$141_3 vdd m1_11381_15778# m1_10560_16202# m1_10299_17343# pfet$141
Xnfet$162_11 m1_22222_21786# m1_22222_21786# vss vss m1_21060_21586# vss nfet$162
Xnfet$157_11 m1_27031_17343# vss m1_27190_17836# vss nfet$157
Xnfet$169_6 m1_1578_16080# m1_1578_16080# vss vss m1_3141_17358# vss nfet$169
Xnfet$176_7 m1_n3822_21786# m1_n3822_21786# m1_n4485_21904# m1_n4485_21904# m1_n3724_21430#
+ vss nfet$176
Xpfet$159_4 vdd m1_28113_15778# m1_27292_16202# m1_27031_17343# pfet$159
Xpfet$141_19 vdd m1_3015_15778# m1_2194_16202# m1_1933_17343# pfet$141
Xpfet$166_5 vdd vdd m1_n4847_25662# m1_n10452_25858# pfet$166
Xnfet$153_9 sd5 vss m1_9331_15478# vss nfet$153
Xnfet$165_0 m1_31535_22102# m1_32818_21586# vss vss nfet$165
Xnfet$154_12 m1_14556_21786# vss m1_15188_21786# vss nfet$154
Xnfet$170_11 m1_15171_20152# m1_15171_20152# m1_n3822_21786# m1_n3822_21786# m1_14005_20470#
+ vss nfet$170
Xnfet$172_1 m1_n6433_17343# m1_n4377_15778# m1_n4994_16080# vss nfet$172
Xpfet$157_1 vdd vdd vdd m1_33050_19550# m1_31535_19792# m1_31535_19792# pfet$157
Xpfet$164_2 vdd m1_n3651_26174# vdd m1_n4978_24224# pfet$164
Xnfet$149_23 m1_25424_24346# m1_25424_24346# m1_24309_25858# m1_24309_25858# m1_26371_25502#
+ vss nfet$149
Xnfet$149_12 m1_17058_24346# m1_17058_24346# m1_15943_25858# m1_15943_25858# m1_18005_25502#
+ vss nfet$149
Xnfet$151_6 m1_2384_21590# m1_2384_21590# m1_3871_22513# m1_3871_22513# m1_2843_21586#
+ vss nfet$151
Xpfet$143_7 vdd vdd vdd m1_6975_19550# m1_965_15478# m1_965_15478# pfet$143
Xnfet$151_13 m1_16452_21590# m1_16452_21590# m1_17939_22513# m1_17939_22513# m1_16911_21586#
+ vss nfet$151
Xpfet$141_4 vdd m1_9485_17714# vdd m1_10560_16202# pfet$141
Xnfet$162_12 m1_18073_21786# m1_18073_21786# vss vss m1_16911_21586# vss nfet$162
Xnfet$157_12 m1_28470_16080# vss m1_28113_15778# vss nfet$157
Xnfet$169_7 m1_5761_16080# m1_5761_16080# m1_5302_17714# m1_5302_17714# m1_5859_16398#
+ vss nfet$169
Xnfet$176_8 m1_9624_19404# m1_9624_19404# vss vss m1_n3724_21430# vss nfet$176
Xpfet$166_6 vdd vdd m1_n4623_25487# fin pfet$166
Xpfet$159_5 vdd m1_29087_15778# m1_28470_16080# m1_27190_17836# pfet$159
Xnfet$154_13 m1_16322_21786# vss m1_16452_21590# vss nfet$154
Xnfet$170_12 m1_18688_20152# m1_18688_20152# m1_n1927_20274# m1_n1927_20274# m1_17522_20470#
+ vss nfet$170
Xnfet$172_2 m1_n6274_17836# m1_n5351_15778# m1_n6172_16202# vss nfet$172
Xpfet$157_2 vdd m1_32818_21586# m1_32818_21586# m1_33050_22344# m1_30256_22102# m1_30256_22102#
+ pfet$157
Xnfet$158_0 m1_n10452_25858# vss m1_n1271_25858# vss nfet$158
Xpfet$164_3 vdd vdd m1_n3651_26174# m1_n3541_23922# pfet$164
Xnfet$149_24 m1_30095_25658# m1_30095_25658# vss vss m1_30554_25502# vss nfet$149
Xnfet$149_13 m1_13363_25658# m1_13363_25658# vss vss m1_13822_25502# vss nfet$149
Xpfet$142_30 vdd vdd vdd m1_17539_22402# m1_16322_21786# m1_16322_21786# pfet$142
Xnfet$151_7 m1_5771_21786# m1_5771_21786# m1_7388_22513# m1_7388_22513# m1_6992_21586#
+ vss nfet$151
Xpfet$143_8 vdd m1_9624_19404# m1_9624_19404# m1_10492_19550# m1_4832_17714# m1_4832_17714#
+ pfet$143
Xpfet$162_0 vdd m1_n10309_25662# m1_n10572_23922# m1_n10796_25662# pfet$162
Xnfet$151_14 m1_12805_21786# m1_12805_21786# m1_14422_22513# m1_14422_22513# m1_14026_21586#
+ vss nfet$151
Xpfet$141_5 vdd m1_7198_15778# m1_6377_16202# m1_6116_17343# pfet$141
Xnfet$162_13 m1_18705_21786# m1_18705_21786# vss vss m1_17543_21586# vss nfet$162
Xnfet$157_13 m1_26217_17714# vss m1_25747_17714# vss nfet$157
Xnfet$169_8 m1_3015_15778# m1_3015_15778# m1_2905_18030# m1_2905_18030# m1_3141_17358#
+ vss nfet$169
Xnfet$176_9 m1_n6380_21786# m1_n6380_21786# m1_n6839_21786# m1_n6839_21786# m1_n6282_21430#
+ vss nfet$176
Xpfet$159_6 vdd m1_28470_16080# m1_28003_18030# m1_27031_17343# pfet$159
Xpfet$166_7 vdd vdd m1_n3541_23922# m1_n3184_24224# pfet$166
Xnfet$154_14 m1_19839_21786# vss m1_19969_21590# vss nfet$154
Xnfet$170_13 m1_13514_15478# m1_13514_15478# m1_n1927_20274# m1_n1927_20274# m1_16890_20470#
+ vss nfet$170
Xnfet$172_3 m1_n6433_17343# m1_n6172_16202# m1_n6657_17518# vss nfet$172
Xnfet$158_1 m1_n789_25858# vss m1_n647_25662# vss nfet$158
Xpfet$164_4 vdd m1_n10452_25858# vdd m1_n4362_24346# pfet$164
Xpfet$142_31 vdd vdd vdd m1_27462_22102# m1_27003_21590# m1_27003_21590# pfet$142
Xnfet$149_14 m1_12875_24346# m1_12875_24346# m1_11760_25858# m1_11760_25858# m1_13822_25502#
+ vss nfet$149
Xpfet$142_20 vdd vdd vdd m1_20428_22102# m1_19969_21590# m1_19969_21590# pfet$142
Xnfet$149_25 m1_29607_24346# m1_29607_24346# m1_28492_25858# m1_28492_25858# m1_30554_25502#
+ vss nfet$149
Xnfet$151_8 m1_23486_21590# m1_23486_21590# m1_24973_22513# m1_24973_22513# m1_23945_21586#
+ vss nfet$151
Xnfet$170_0 m1_4620_20152# m1_4620_20152# m1_2590_19404# m1_2590_19404# m1_3454_20470#
+ vss nfet$170
Xpfet$143_9 vdd m1_9624_19404# m1_9624_19404# m1_9856_19850# m1_9418_19550# m1_9418_19550#
+ pfet$143
Xpfet$155_0 vdd vdd vdd m1_36073_22344# define define pfet$155
Xpfet$162_1 vdd m1_n9952_24224# m1_n8848_25658# m1_n10933_25858# pfet$162
Xnfet$151_15 m1_26873_21786# m1_26873_21786# m1_28490_22513# m1_28490_22513# m1_28094_21586#
+ vss nfet$151
Xpfet$141_6 vdd vdd m1_7198_15778# m1_7555_16080# pfet$141
Xnfet$162_14 m1_15188_21786# m1_15188_21786# vss vss m1_14026_21586# vss nfet$162
.ends

.subckt asc_drive_buffer$1 vss in vdd out
Xpfet$208_0 vdd vdd m1_4002_n1060# m1_3466_n454# pfet$208
Xpfet$206_0 out out m1_4274_n1060# vdd m1_4274_n1060# out vdd vdd m1_4274_n1060# out
+ m1_4274_n1060# m1_4274_n1060# out m1_4274_n1060# vdd m1_4274_n1060# vdd m1_4274_n1060#
+ pfet$206
Xnfet$221_0 m1_3466_n454# vss m1_4002_n1060# vss nfet$221
Xnfet$219_0 m1_4274_n1060# vss m1_4002_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ m1_4274_n1060# vss m1_4002_n1060# vss nfet$219
Xpfet$209_0 vdd vdd m1_3466_n454# in pfet$209
Xpfet$207_0 m1_4274_n1060# vdd vdd m1_4274_n1060# m1_4002_n1060# m1_4002_n1060# m1_4274_n1060#
+ vdd m1_4002_n1060# m1_4002_n1060# pfet$207
Xnfet$222_0 in vss m1_3466_n454# vss nfet$222
Xnfet$220_0 out out vss m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# m1_4274_n1060#
+ m1_4274_n1060# out m1_4274_n1060# m1_4274_n1060# out vss m1_4274_n1060# vss vss
+ nfet$220
.ends

.subckt xp_3_1_MUX S0 S1 VDD VSS OUT_1 C_1 B_1 A_1
Xnfet$213_0 S1 VSS m1_n432_n1290# VSS nfet$213
Xnfet$213_1 S0 VSS m1_n432_458# VSS nfet$213
Xpfet$199_0 VDD A_1 m1_239_n318# m1_n432_458# pfet$199
Xpfet$199_1 VDD C_1 OUT_1 S1 pfet$199
Xpfet$199_2 VDD B_1 m1_239_n318# S0 pfet$199
Xpfet$199_3 VDD m1_239_n318# OUT_1 m1_n432_n1290# pfet$199
Xnfet$212_0 m1_n432_n1290# C_1 OUT_1 VSS nfet$212
Xnfet$212_1 m1_n432_458# B_1 m1_239_n318# VSS nfet$212
Xnfet$212_2 S1 m1_239_n318# OUT_1 VSS nfet$212
Xnfet$212_3 S0 A_1 m1_239_n318# VSS nfet$212
Xpfet$200_0 VDD VDD m1_n432_n1290# S1 pfet$200
Xpfet$200_1 VDD VDD m1_n432_458# S0 pfet$200
.ends

.subckt pfet$176 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$189 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pass1u05u$1 VDD VSS ind ins clkn clkp
Xpfet$176_0 VDD ind ins clkp pfet$176
Xnfet$189_0 clkn ind ins VSS nfet$189
.ends

.subckt nfet$188 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt nfet$187 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$173 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_954_0# w_n180_n88# a_854_n136#
+ a_n92_0# a_446_n136# a_650_n136# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt pfet$178 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=0.5u
.ends

.subckt pfet$177 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$190 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt inv1u05u$1 VDD VSS out in
Xpfet$177_0 VDD VDD out in pfet$177
Xnfet$190_0 in VSS out VSS nfet$190
.ends

.subckt nfet$186 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=4.27p pd=15.22u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.82p pd=7.52u as=4.27p ps=15.22u w=7u l=0.5u
.ends

.subckt pfet$175 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=4.55p ps=15.3u w=7u l=0.5u
.ends

.subckt nfet$191 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$174 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_954_0# w_n180_n88#
+ a_38_n60# a_n92_0# a_1058_n60# a_854_n60# a_342_0# a_138_0# a_650_n60#
X0 a_954_0# a_854_n60# a_750_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X1 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X2 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
X3 a_1158_0# a_1058_n60# a_954_0# w_n180_n88# pfet_03v3 ad=4.55p pd=15.3u as=1.82p ps=7.52u w=7u l=0.5u
X4 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=4.55p ps=15.3u w=7u l=0.5u
X5 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=1.82p pd=7.52u as=1.82p ps=7.52u w=7u l=0.5u
.ends

.subckt xp_programmable_basic_pump up vdd s1 s2 s3 s4 down out iref vss
Xpass1u05u$1_2 vdd vss iref pass1u05u$1_2/ins s1 inv1u05u$1_3/out pass1u05u$1
Xnfet$188_1 m1_n7879_n12170# pass1u05u$1_0/ins m1_n7879_n12170# out pass1u05u$1_0/ins
+ vss nfet$188
Xnfet$187_11 vss vss vss vss vss vss nfet$187
Xpfet$173_9 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$173
Xpass1u05u$1_3 vdd vss pass1u05u$1_7/ind pass1u05u$1_3/ins s1 inv1u05u$1_3/out pass1u05u$1
Xnfet$187_12 vss vss vss vss vss vss nfet$187
Xnfet$188_2 vss down vss m1_n7879_n12170# down vss nfet$188
Xpfet$178_0 vdd s3 pass1u05u$1_5/ins vdd pfet$178
Xinv1u05u$1_0 vdd vss inv1u05u$1_0/out s4 inv1u05u$1
Xpass1u05u$1_4 vdd vss pass1u05u$1_7/ind pass1u05u$1_4/ins s2 inv1u05u$1_2/out pass1u05u$1
Xnfet$188_3 vss down vss m1_n7879_n12170# down vss nfet$188
Xnfet$187_13 vss vss vss vss vss vss nfet$187
Xpfet$178_1 vdd s2 pass1u05u$1_4/ins vdd pfet$178
Xnfet$186_0 pass1u05u$1_6/ins pass1u05u$1_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$186
Xinv1u05u$1_1 vdd vss inv1u05u$1_1/out s3 inv1u05u$1
Xpass1u05u$1_5 vdd vss pass1u05u$1_7/ind pass1u05u$1_5/ins s3 inv1u05u$1_1/out pass1u05u$1
Xpfet$175_20 vdd vdd vdd vdd pfet$175
Xnfet$188_4 vss down vss m1_n7879_n12170# down vss nfet$188
Xpfet$178_2 vdd s1 pass1u05u$1_3/ins vdd pfet$178
Xnfet$186_1 pass1u05u$1_6/ins pass1u05u$1_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$186
Xinv1u05u$1_2 vdd vss inv1u05u$1_2/out s2 inv1u05u$1
Xpfet$175_21 vdd vdd vdd vdd pfet$175
Xpass1u05u$1_6 vdd vss iref pass1u05u$1_6/ins s4 inv1u05u$1_0/out pass1u05u$1
Xnfet$188_5 vss down vss m1_n7879_n12170# down vss nfet$188
Xpfet$175_10 vdd vdd vdd vdd pfet$175
Xpfet$178_3 vdd s4 pass1u05u$1_7/ins vdd pfet$178
Xnfet$186_2 pass1u05u$1_6/ins pass1u05u$1_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$186
Xnfet$191_0 inv1u05u$1_2/out pass1u05u$1_1/ins vss vss nfet$191
Xinv1u05u$1_3 vdd vss inv1u05u$1_3/out s1 inv1u05u$1
Xpass1u05u$1_7 vdd vss pass1u05u$1_7/ind pass1u05u$1_7/ins s4 inv1u05u$1_0/out pass1u05u$1
Xpfet$175_22 vdd vdd vdd vdd pfet$175
Xnfet$188_6 m1_n7879_n12170# pass1u05u$1_0/ins m1_n7879_n12170# out pass1u05u$1_0/ins
+ vss nfet$188
Xpfet$175_11 vdd vdd vdd vdd pfet$175
Xnfet$191_1 inv1u05u$1_3/out pass1u05u$1_2/ins vss vss nfet$191
Xnfet$186_3 vss vss vss vss vss vss nfet$186
Xpfet$175_23 vdd vdd vdd vdd pfet$175
Xnfet$188_7 m1_n7879_n12170# pass1u05u$1_0/ins m1_n7879_n12170# out pass1u05u$1_0/ins
+ vss nfet$188
Xpfet$175_12 vdd vdd vdd vdd pfet$175
Xnfet$186_4 pass1u05u$1_6/ins pass1u05u$1_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$186
Xnfet$191_2 inv1u05u$1_0/out pass1u05u$1_6/ins vss vss nfet$191
Xpfet$175_13 vdd vdd vdd vdd pfet$175
Xnfet$188_8 vss vdd vss m1_n8144_n9165# vdd vss nfet$188
Xnfet$191_3 inv1u05u$1_1/out pass1u05u$1_0/ins vss vss nfet$191
Xnfet$186_5 vss vss vss vss vss vss nfet$186
Xpfet$174_0 vdd vdd m1_n4127_3649# vss vss m1_n4127_3649# vdd vss vdd vss vss vdd
+ m1_n4127_3649# vss pfet$174
Xpfet$175_14 vdd vdd vdd vdd pfet$175
Xnfet$186_6 pass1u05u$1_6/ins pass1u05u$1_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$186
Xnfet$188_9 m1_n7216_n8262# iref m1_n7216_n8262# pass1u05u$1_7/ind iref vss nfet$188
Xpfet$174_1 m1_n5580_883# m1_n5580_883# out pass1u05u$1_5/ins pass1u05u$1_5/ins out
+ vdd pass1u05u$1_5/ins m1_n5580_883# pass1u05u$1_5/ins pass1u05u$1_5/ins m1_n5580_883#
+ out pass1u05u$1_5/ins pfet$174
Xpfet$175_15 vdd vdd vdd vdd pfet$175
Xnfet$186_7 pass1u05u$1_6/ins pass1u05u$1_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$186
Xpfet$174_2 m1_n5580_883# m1_n5580_883# out pass1u05u$1_5/ins pass1u05u$1_5/ins out
+ vdd pass1u05u$1_5/ins m1_n5580_883# pass1u05u$1_5/ins pass1u05u$1_5/ins m1_n5580_883#
+ out pass1u05u$1_5/ins pfet$174
Xpfet$175_16 vdd vdd vdd vdd pfet$175
Xnfet$186_8 pass1u05u$1_6/ins pass1u05u$1_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$186
Xpfet$174_3 m1_n5580_883# m1_n5580_883# out pass1u05u$1_5/ins pass1u05u$1_5/ins out
+ vdd pass1u05u$1_5/ins m1_n5580_883# pass1u05u$1_5/ins pass1u05u$1_5/ins m1_n5580_883#
+ out pass1u05u$1_5/ins pfet$174
Xpfet$175_17 vdd vdd vdd vdd pfet$175
Xnfet$188_10 m1_n8607_n8040# pass1u05u$1_1/ins m1_n8607_n8040# out pass1u05u$1_1/ins
+ vss nfet$188
Xnfet$186_9 pass1u05u$1_6/ins pass1u05u$1_6/ins m1_n8807_n11192# m1_n8807_n11192#
+ out vss nfet$186
Xpfet$174_4 m1_n5580_883# m1_n5580_883# out pass1u05u$1_5/ins pass1u05u$1_5/ins out
+ vdd pass1u05u$1_5/ins m1_n5580_883# pass1u05u$1_5/ins pass1u05u$1_5/ins m1_n5580_883#
+ out pass1u05u$1_5/ins pfet$174
Xpfet$175_18 vdd vdd vdd vdd pfet$175
Xnfet$188_11 m1_n8144_n9165# iref m1_n8144_n9165# iref iref vss nfet$188
Xpfet$174_5 m1_n4127_3649# m1_n4127_3649# pass1u05u$1_7/ind pass1u05u$1_7/ind pass1u05u$1_7/ind
+ pass1u05u$1_7/ind vdd pass1u05u$1_7/ind m1_n4127_3649# pass1u05u$1_7/ind pass1u05u$1_7/ind
+ m1_n4127_3649# pass1u05u$1_7/ind pass1u05u$1_7/ind pfet$174
Xpfet$175_19 vdd vdd vdd vdd pfet$175
Xnfet$188_12 vss down vss m1_n8607_n8040# down vss nfet$188
Xnfet$188_13 vss vdd vss m1_n7216_n8262# vdd vss nfet$188
Xpfet$173_20 m1_n8156_628# m1_n8156_628# pass1u05u$1_7/ins out out vdd pass1u05u$1_7/ins
+ m1_n8156_628# pass1u05u$1_7/ins pass1u05u$1_7/ins m1_n8156_628# out pass1u05u$1_7/ins
+ pass1u05u$1_7/ins pfet$173
Xnfet$188_14 m1_n8607_n8040# pass1u05u$1_1/ins m1_n8607_n8040# out pass1u05u$1_1/ins
+ vss nfet$188
Xpfet$173_21 m1_n6703_2564# m1_n6703_2564# pass1u05u$1_4/ins out out vdd pass1u05u$1_4/ins
+ m1_n6703_2564# pass1u05u$1_4/ins pass1u05u$1_4/ins m1_n6703_2564# out pass1u05u$1_4/ins
+ pass1u05u$1_4/ins pfet$173
Xpfet$173_10 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$173
Xnfet$188_15 vss down vss m1_n8607_n8040# down vss nfet$188
Xpfet$173_22 m1_n8156_628# m1_n8156_628# pass1u05u$1_7/ins out out vdd pass1u05u$1_7/ins
+ m1_n8156_628# pass1u05u$1_7/ins pass1u05u$1_7/ins m1_n8156_628# out pass1u05u$1_7/ins
+ pass1u05u$1_7/ins pfet$173
Xpfet$173_11 vdd vdd up m1_n5450_4559# m1_n5450_4559# vdd up vdd up up vdd m1_n5450_4559#
+ up up pfet$173
Xpfet$173_23 m1_n8156_628# m1_n8156_628# pass1u05u$1_7/ins out out vdd pass1u05u$1_7/ins
+ m1_n8156_628# pass1u05u$1_7/ins pass1u05u$1_7/ins m1_n8156_628# out pass1u05u$1_7/ins
+ pass1u05u$1_7/ins pfet$173
Xpfet$173_12 vdd vdd up m1_n6703_2564# m1_n6703_2564# vdd up vdd up up vdd m1_n6703_2564#
+ up up pfet$173
Xpfet$173_24 m1_n5450_4559# m1_n5450_4559# pass1u05u$1_3/ins out out vdd pass1u05u$1_3/ins
+ m1_n5450_4559# pass1u05u$1_3/ins pass1u05u$1_3/ins m1_n5450_4559# out pass1u05u$1_3/ins
+ pass1u05u$1_3/ins pfet$173
Xnfet$187_0 down down vss vss m1_n8807_n11192# vss nfet$187
Xpfet$173_13 vdd vdd up m1_n6703_2564# m1_n6703_2564# vdd up vdd up up vdd m1_n6703_2564#
+ up up pfet$173
Xpfet$173_25 m1_n6703_2564# m1_n6703_2564# pass1u05u$1_4/ins out out vdd pass1u05u$1_4/ins
+ m1_n6703_2564# pass1u05u$1_4/ins pass1u05u$1_4/ins m1_n6703_2564# out pass1u05u$1_4/ins
+ pass1u05u$1_4/ins pfet$173
Xpfet$173_14 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$173
Xnfet$187_1 down down vss vss m1_n8807_n11192# vss nfet$187
Xnfet$187_2 down down vss vss m1_n8807_n11192# vss nfet$187
Xpfet$173_15 m1_n8156_628# m1_n8156_628# pass1u05u$1_7/ins out out vdd pass1u05u$1_7/ins
+ m1_n8156_628# pass1u05u$1_7/ins pass1u05u$1_7/ins m1_n8156_628# out pass1u05u$1_7/ins
+ pass1u05u$1_7/ins pfet$173
Xnfet$187_3 down down vss vss m1_n8807_n11192# vss nfet$187
Xpfet$173_16 m1_n8156_628# m1_n8156_628# pass1u05u$1_7/ins out out vdd pass1u05u$1_7/ins
+ m1_n8156_628# pass1u05u$1_7/ins pass1u05u$1_7/ins m1_n8156_628# out pass1u05u$1_7/ins
+ pass1u05u$1_7/ins pfet$173
Xpfet$173_17 m1_n8156_628# m1_n8156_628# pass1u05u$1_7/ins out out vdd pass1u05u$1_7/ins
+ m1_n8156_628# pass1u05u$1_7/ins pass1u05u$1_7/ins m1_n8156_628# out pass1u05u$1_7/ins
+ pass1u05u$1_7/ins pfet$173
Xnfet$187_4 vss vss vss vss vss vss nfet$187
Xnfet$186_10 pass1u05u$1_2/ins pass1u05u$1_2/ins m1_n7679_n8960# m1_n7679_n8960# out
+ vss nfet$186
Xpfet$173_18 m1_n8156_628# m1_n8156_628# pass1u05u$1_7/ins out out vdd pass1u05u$1_7/ins
+ m1_n8156_628# pass1u05u$1_7/ins pass1u05u$1_7/ins m1_n8156_628# out pass1u05u$1_7/ins
+ pass1u05u$1_7/ins pfet$173
Xnfet$187_5 vss vss vss vss vss vss nfet$187
Xnfet$186_11 vss vss vss vss vss vss nfet$186
Xpfet$175_0 vdd vdd vdd vdd pfet$175
Xpfet$173_19 m1_n8156_628# m1_n8156_628# pass1u05u$1_7/ins out out vdd pass1u05u$1_7/ins
+ m1_n8156_628# pass1u05u$1_7/ins pass1u05u$1_7/ins m1_n8156_628# out pass1u05u$1_7/ins
+ pass1u05u$1_7/ins pfet$173
Xnfet$187_6 down down vss vss m1_n8807_n11192# vss nfet$187
Xnfet$186_12 down down vss vss m1_n7679_n8960# vss nfet$186
Xpfet$175_1 vdd vdd vdd vdd pfet$175
Xnfet$186_13 vss vss vss vss vss vss nfet$186
Xnfet$187_7 down down vss vss m1_n8807_n11192# vss nfet$187
Xpfet$175_2 vdd vdd vdd vdd pfet$175
Xnfet$186_14 vss vss vss vss vss vss nfet$186
Xnfet$187_8 down down vss vss m1_n8807_n11192# vss nfet$187
Xpfet$175_3 vdd vdd vdd vdd pfet$175
Xpfet$173_0 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$173
Xnfet$186_15 vss vss vss vss vss vss nfet$186
Xnfet$187_9 down down vss vss m1_n8807_n11192# vss nfet$187
Xpfet$173_1 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$173
Xpfet$175_4 vdd vdd vdd vdd pfet$175
Xpfet$175_5 vdd vdd vdd vdd pfet$175
Xpfet$173_2 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$173
Xpfet$175_6 vdd vdd vdd vdd pfet$175
Xpfet$173_3 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$173
Xpfet$175_7 vdd vdd vdd vdd pfet$175
Xpfet$173_4 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$173
Xpfet$175_8 vdd vdd vdd vdd pfet$175
Xpfet$173_5 vdd vdd up m1_n5580_883# m1_n5580_883# vdd up vdd up up vdd m1_n5580_883#
+ up up pfet$173
Xpfet$173_6 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$173
Xpfet$175_9 vdd vdd vdd vdd pfet$175
Xpass1u05u$1_0 vdd vss iref pass1u05u$1_0/ins s3 inv1u05u$1_1/out pass1u05u$1
Xpfet$173_7 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$173
Xpass1u05u$1_1 vdd vss iref pass1u05u$1_1/ins s2 inv1u05u$1_2/out pass1u05u$1
Xnfet$187_10 vss vss vss vss vss vss nfet$187
Xnfet$188_0 m1_n7879_n12170# pass1u05u$1_0/ins m1_n7879_n12170# out pass1u05u$1_0/ins
+ vss nfet$188
Xpfet$173_8 vdd vdd up m1_n8156_628# m1_n8156_628# vdd up vdd up up vdd m1_n8156_628#
+ up up pfet$173
.ends

.subckt asc_hysteresis_buffer$1 vss in vdd out
Xnfet$193_0 m1_348_648# vss m1_884_42# vss nfet$193
Xpfet$183_0 vdd vdd m1_884_42# m1_1156_42# pfet$183
Xpfet$181_0 vdd vdd m1_348_648# in pfet$181
Xnfet$196_0 m1_1156_42# vss m1_884_42# vss nfet$196
Xpfet$179_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd
+ m1_884_42# m1_884_42# pfet$179
Xnfet$194_0 in vss m1_348_648# vss nfet$194
Xnfet$192_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$192
Xpfet$182_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$182
Xpfet$180_0 vdd vdd m1_884_42# m1_348_648# pfet$180
Xnfet$195_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$195
.ends

.subckt pfet$219 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$212 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$210 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$236 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$229 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$234 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt nfet$227 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$232 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$217 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$225 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$222 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$230 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$215 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt nfet$223 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$220 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt pfet$213 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$211 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$235 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt nfet$228 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt nfet$233 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$218 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt nfet$226 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$231 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt pfet$216 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$224 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$221 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt pfet$214 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt asc_PFD_DFF_20250831 vss down up vdd fref fdiv
Xpfet$219_10 vdd vdd m1_3349_n9089# m1_2779_n10883# pfet$219
Xpfet$212_2 vdd vdd m1_2068_n5361# m1_2758_n8889# pfet$212
Xpfet$219_11 vdd vdd down m1_2779_n10883# pfet$219
Xpfet$212_3 vdd vdd m1_1452_n5483# m1_832_n5785# pfet$212
Xpfet$210_0 vdd m1_832_n5785# m1_1096_n5165# m1_n3885_n6084# pfet$210
Xnfet$236_0 up up m1_5895_n8089# m1_5895_n8089# m1_5043_n9245# vss nfet$236
Xpfet$219_12 vdd m1_2556_n10129# m1_3349_n9089# m1_n3884_n11124# pfet$219
Xpfet$212_4 vdd vdd m1_1095_n4045# vdd pfet$212
Xpfet$210_1 vdd m1_1452_n5483# m1_2556_n4049# m1_n3885_n6084# pfet$210
Xnfet$236_1 down down vss vss m1_5043_n9245# vss nfet$236
Xpfet$219_13 vdd vdd m1_n5427_n8573# m1_n4677_n8889# pfet$219
Xnfet$229_0 m1_n5428_n3533# vss m1_n3885_n4045# vss nfet$229
Xpfet$210_2 vdd m1_1095_n4045# m1_832_n5785# m1_n3885_n4045# pfet$210
Xpfet$219_14 vdd vdd m1_n3884_n11124# m1_n5427_n10882# pfet$219
Xnfet$229_1 m1_n5868_n3849# vss m1_n5650_n4045# vss nfet$229
Xpfet$210_3 vdd m1_2556_n4049# m1_3349_n5165# m1_n3885_n4045# pfet$210
Xpfet$219_15 vdd m1_n5427_n10882# vdd m1_n5649_n11124# pfet$219
Xnfet$229_2 m1_n5428_n5842# vss m1_n3885_n6084# vss nfet$229
Xpfet$219_0 vdd vdd m1_2779_n10883# m1_2068_n8889# pfet$219
Xnfet$234_0 m1_n3884_n11124# vss m1_n3098_n10720# vss nfet$234
Xpfet$219_16 vdd vdd m1_n5427_n10882# m1_n4677_n10522# pfet$219
Xpfet$219_1 vdd m1_2779_n10883# vdd m1_2556_n10129# pfet$219
Xnfet$234_1 m1_n3884_n9085# vss m1_n3098_n9135# vss nfet$234
Xnfet$229_3 fref vss m1_n5868_n3849# vss nfet$229
Xnfet$227_0 m1_5895_n8089# vss m1_5464_n5483# vss nfet$227
Xpfet$219_17 vdd vdd m1_n5649_n11124# m1_n5867_n10544# pfet$219
Xpfet$219_2 vdd m1_1095_n11125# m1_832_n8573# m1_n3884_n11124# pfet$219
Xnfet$227_1 m1_5464_n5483# vss m1_4978_n5483# vss nfet$227
Xpfet$219_18 vdd vdd m1_n5867_n10544# fdiv pfet$219
Xnfet$232_0 m1_2556_n10129# m1_2556_n10129# vss vss m1_3015_n10205# vss nfet$232
Xpfet$219_3 vdd m1_1452_n8889# m1_2556_n10129# m1_n3884_n9085# pfet$219
Xpfet$217_0 vdd m1_n5428_n3533# vdd m1_n5650_n4045# pfet$217
Xpfet$219_19 vdd vdd m1_n3884_n9085# m1_n5427_n8573# pfet$219
Xpfet$219_4 vdd vdd m1_1452_n8889# m1_832_n8573# pfet$219
Xnfet$232_1 m1_1452_n8889# m1_1452_n8889# m1_1096_n9089# m1_1096_n9089# m1_1550_n9245#
+ vss nfet$232
Xpfet$217_1 vdd vdd m1_n5428_n3533# m1_n4678_n3849# pfet$217
Xnfet$225_0 m1_2779_n3533# vss up vss nfet$225
Xpfet$219_5 vdd vdd m1_1095_n11125# vdd pfet$219
Xnfet$232_2 m1_2068_n8889# m1_2068_n8889# vss vss m1_1550_n9245# vss nfet$232
Xpfet$217_2 vdd m1_n5428_n5842# vdd m1_n5868_n3849# pfet$217
Xnfet$225_1 m1_2779_n3533# vss m1_3349_n5165# vss nfet$225
Xpfet$222_0 vdd m1_5895_n8089# vdd down pfet$222
Xpfet$219_6 vdd vdd m1_1096_n9089# m1_1452_n8889# pfet$219
Xnfet$225_2 m1_2758_n8889# vss m1_2068_n5361# vss nfet$225
Xpfet$222_1 vdd vdd m1_5895_n8089# up pfet$222
Xnfet$232_3 m1_2068_n8889# m1_2068_n8889# m1_2779_n10883# m1_2779_n10883# m1_3015_n10205#
+ vss nfet$232
Xnfet$230_0 m1_n4678_n3849# m1_n4678_n3849# m1_n5428_n3533# m1_n5428_n3533# m1_n5192_n4205#
+ vss nfet$230
Xpfet$217_3 vdd vdd m1_n5428_n5842# m1_n4678_n5482# pfet$217
Xpfet$215_0 m1_n1926_n4095# vdd vdd m1_n3099_n4095# pfet$215
Xnfet$225_3 m1_832_n5785# vss m1_1452_n5483# vss nfet$225
Xpfet$219_7 vdd m1_832_n8573# m1_1096_n9089# m1_n3884_n9085# pfet$219
Xnfet$232_4 m1_n4677_n10522# m1_n4677_n10522# m1_n5427_n10882# m1_n5427_n10882# m1_n5191_n10204#
+ vss nfet$232
Xnfet$223_0 m1_n3885_n4045# m1_832_n5785# m1_1096_n5165# vss nfet$223
Xpfet$215_1 m1_n4678_n3849# vdd vdd m1_n1926_n5680# pfet$215
Xnfet$230_1 m1_n5650_n4045# m1_n5650_n4045# vss vss m1_n5192_n4205# vss nfet$230
Xpfet$219_8 vdd m1_1096_n9089# vdd m1_2068_n8889# pfet$219
Xnfet$225_4 vdd vss m1_1095_n4045# vss nfet$225
Xnfet$223_1 m1_n3885_n4045# m1_1452_n5483# m1_2556_n4049# vss nfet$223
Xnfet$232_5 m1_n5649_n11124# m1_n5649_n11124# vss vss m1_n5191_n10204# vss nfet$232
Xnfet$230_2 m1_n4678_n5482# m1_n4678_n5482# m1_n5428_n5842# m1_n5428_n5842# m1_n5192_n5164#
+ vss nfet$230
Xpfet$220_0 vdd vdd m1_n3098_n10720# m1_n3884_n11124# pfet$220
Xpfet$215_2 m1_n1926_n5680# vdd vdd m1_n3099_n5680# pfet$215
Xpfet$219_9 vdd vdd m1_2068_n8889# m1_2758_n8889# pfet$219
Xnfet$232_6 m1_n4677_n8889# m1_n4677_n8889# m1_n5427_n8573# m1_n5427_n8573# m1_n5191_n9245#
+ vss nfet$232
Xnfet$223_2 m1_n3885_n6084# m1_1095_n4045# m1_832_n5785# vss nfet$223
Xnfet$230_3 m1_n5868_n3849# m1_n5868_n3849# vss vss m1_n5192_n5164# vss nfet$230
Xpfet$215_3 m1_n4678_n5482# vdd vdd m1_n1926_n4095# pfet$215
Xpfet$220_1 vdd vdd m1_n3098_n9135# m1_n3884_n9085# pfet$220
Xpfet$213_0 vdd vdd m1_2758_n8889# m1_4978_n5483# pfet$213
Xnfet$232_7 m1_n5867_n10544# m1_n5867_n10544# vss vss m1_n5191_n9245# vss nfet$232
Xnfet$223_3 m1_n3885_n6084# m1_2556_n4049# m1_3349_n5165# vss nfet$223
Xpfet$211_0 vdd vdd m1_1096_n5165# m1_1452_n5483# pfet$211
Xpfet$211_1 vdd m1_1096_n5165# vdd m1_2068_n5361# pfet$211
Xpfet$211_2 vdd m1_2779_n3533# vdd m1_2556_n4049# pfet$211
Xpfet$211_3 vdd vdd m1_2779_n3533# m1_2068_n5361# pfet$211
Xnfet$235_0 m1_n4677_n8889# m1_n1925_n10720# vss vss nfet$235
Xnfet$235_1 m1_n1925_n10720# m1_n3098_n10720# vss vss nfet$235
Xnfet$228_0 m1_n1926_n4095# m1_n3099_n4095# vss vss nfet$228
Xnfet$235_2 m1_n4677_n10522# m1_n1925_n9135# vss vss nfet$235
Xnfet$228_1 m1_n4678_n3849# m1_n1926_n5680# vss vss nfet$228
Xnfet$233_0 m1_n3884_n9085# m1_1095_n11125# m1_832_n8573# vss nfet$233
Xnfet$235_3 m1_n1925_n9135# m1_n3098_n9135# vss vss nfet$235
Xnfet$228_2 m1_n1926_n5680# m1_n3099_n5680# vss vss nfet$228
Xpfet$218_0 vdd vdd m1_n3099_n4095# m1_n3885_n4045# pfet$218
Xnfet$228_3 m1_n4678_n5482# m1_n1926_n4095# vss vss nfet$228
Xnfet$233_1 m1_n3884_n11124# m1_1452_n8889# m1_2556_n10129# vss nfet$233
Xpfet$218_1 vdd vdd m1_n3099_n5680# m1_n3885_n6084# pfet$218
Xnfet$226_0 m1_4978_n5483# vss m1_2758_n8889# vss nfet$226
Xnfet$233_2 m1_832_n8573# vss m1_1452_n8889# vss nfet$233
Xnfet$233_3 vdd vss m1_1095_n11125# vss nfet$233
Xnfet$231_0 m1_n3885_n4045# vss m1_n3099_n4095# vss nfet$231
Xpfet$216_0 vdd vdd m1_n3885_n4045# m1_n5428_n3533# pfet$216
Xnfet$224_0 m1_2068_n5361# m1_2068_n5361# vss vss m1_1550_n5165# vss nfet$224
Xnfet$233_4 m1_n3884_n11124# m1_832_n8573# m1_1096_n9089# vss nfet$233
Xnfet$231_1 m1_n3885_n6084# vss m1_n3099_n5680# vss nfet$231
Xpfet$216_1 vdd vdd m1_n5650_n4045# m1_n5868_n3849# pfet$216
Xnfet$233_5 m1_2758_n8889# vss m1_2068_n8889# vss nfet$233
Xnfet$224_1 m1_1452_n5483# m1_1452_n5483# m1_1096_n5165# m1_1096_n5165# m1_1550_n5165#
+ vss nfet$224
Xnfet$233_10 m1_n5867_n10544# vss m1_n5649_n11124# vss nfet$233
Xpfet$216_2 vdd vdd m1_n3885_n6084# m1_n5428_n5842# pfet$216
Xpfet$221_0 m1_n4677_n8889# vdd vdd m1_n1925_n10720# pfet$221
Xnfet$224_2 m1_2556_n4049# m1_2556_n4049# vss vss m1_3015_n4205# vss nfet$224
Xnfet$233_6 m1_2779_n10883# vss down vss nfet$233
Xnfet$233_11 fdiv vss m1_n5867_n10544# vss nfet$233
Xpfet$221_1 m1_n1925_n10720# vdd vdd m1_n3098_n10720# pfet$221
Xpfet$216_3 vdd vdd m1_n5868_n3849# fref pfet$216
Xpfet$214_0 vdd vdd m1_5464_n5483# m1_5895_n8089# pfet$214
Xnfet$233_7 m1_2779_n10883# vss m1_3349_n9089# vss nfet$233
Xnfet$224_3 m1_2068_n5361# m1_2068_n5361# m1_2779_n3533# m1_2779_n3533# m1_3015_n4205#
+ vss nfet$224
Xnfet$233_12 m1_n5427_n8573# vss m1_n3884_n9085# vss nfet$233
Xpfet$221_2 m1_n4677_n10522# vdd vdd m1_n1925_n9135# pfet$221
Xpfet$214_1 vdd vdd m1_4978_n5483# m1_5464_n5483# pfet$214
Xnfet$233_8 m1_n3884_n9085# m1_2556_n10129# m1_3349_n9089# vss nfet$233
Xpfet$221_3 m1_n1925_n9135# vdd vdd m1_n3098_n9135# pfet$221
Xnfet$233_9 m1_n5427_n10882# vss m1_n3884_n11124# vss nfet$233
Xpfet$212_0 vdd vdd m1_3349_n5165# m1_2779_n3533# pfet$212
Xpfet$219_20 vdd m1_n5427_n8573# vdd m1_n5867_n10544# pfet$219
Xpfet$212_1 vdd vdd up m1_2779_n3533# pfet$212
.ends

.subckt pfet$223 a_254_0# a_348_560# w_n180_n88# a_414_0# a_n92_0# a_94_0# a_574_0#
+ a_508_560# a_188_560# a_28_560#
X0 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$237 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt BIAS vdd vss 100n 200n res 200p1 200p2
Xpfet$223_9 vdd res vdd 100n vdd 100n vdd res res res pfet$223
Xnfet$237_0 m1_27_n1423# vss 200p1 m1_27_n1423# vss 200p1 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$237
Xnfet$237_1 vss vss vss vss vss vss vss vss vss vss nfet$237
Xnfet$237_2 m1_27_n1423# vss 200p2 m1_27_n1423# vss 200p2 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$237
Xnfet$237_3 vss vss vss vss vss vss vss vss vss vss nfet$237
Xnfet$237_5 m1_27_n1423# vss 200p1 m1_27_n1423# vss 200p1 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$237
Xnfet$237_4 m1_27_n1423# vss 200p2 m1_27_n1423# vss 200p2 m1_27_n1423# vss m1_27_n1423#
+ vss nfet$237
Xpfet$223_10 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$223
Xnfet$237_6 m1_27_n1423# vss m1_27_n1423# m1_27_n1423# vss m1_27_n1423# m1_27_n1423#
+ vss m1_27_n1423# vss nfet$237
Xpfet$223_12 vdd res vdd 100n vdd 100n vdd res res res pfet$223
Xpfet$223_11 vdd res vdd 200n vdd 200n vdd res res res pfet$223
Xnfet$237_7 m1_27_n1423# vss m1_27_n1423# m1_27_n1423# vss m1_27_n1423# m1_27_n1423#
+ vss m1_27_n1423# vss nfet$237
Xpfet$223_13 vdd res vdd res vdd res vdd res res res pfet$223
Xpfet$223_14 vdd res vdd 200n vdd 200n vdd res res res pfet$223
Xpfet$223_0 vdd res vdd 200n vdd 200n vdd res res res pfet$223
Xpfet$223_15 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$223
Xpfet$223_2 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$223
Xpfet$223_1 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$223
Xpfet$223_3 vdd res vdd m1_27_n1423# vdd m1_27_n1423# vdd res res res pfet$223
Xpfet$223_4 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$223
Xpfet$223_5 vdd res vdd 200n vdd 200n vdd res res res pfet$223
Xpfet$223_6 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$223
Xpfet$223_7 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$223
Xpfet$223_8 vdd res vdd res vdd res vdd res res res pfet$223
.ends

.subckt pfet$224 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=9.75p pd=31.3u as=9.75p ps=31.3u w=15u l=0.5u
.ends

.subckt nfet$238 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.5u
.ends

.subckt pfet$226 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt cap_mim$4 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=10u c_length=5u
.ends

.subckt nfet$239 a_n84_0# a_38_n132# a_138_0# VSUBS
X0 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=3.05p pd=11.22u as=3.05p ps=11.22u w=5u l=0.5u
.ends

.subckt pfet$225 w_n180_n88# a_38_n60# a_n92_0# a_138_0#
X0 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=9.75p pd=31.3u as=9.75p ps=31.3u w=15u l=0.5u
.ends

.subckt nfet$240 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt CSRVCO_20250823 vctrl vosc vdd vss
Xpfet$224_11 vdd m1_n12264_2422# m1_n11916_1270# m1_n9352_266# pfet$224
Xpfet$224_10 vdd m1_n14208_3657# m1_n10810_266# m1_n11296_266# pfet$224
Xnfet$238_1 vctrl vss m1_n12268_985# vss nfet$238
Xnfet$238_2 vctrl vss m1_n14283_186# vss nfet$238
Xpfet$224_12 vdd m1_n14693_3963# m1_n11296_266# m1_n11782_266# pfet$224
Xnfet$238_3 vctrl vss m1_n13794_186# vss nfet$238
Xpfet$224_13 vdd m1_n13722_3340# m1_n10324_266# m1_n10810_266# pfet$224
Xnfet$238_4 vctrl vss m1_n13240_368# vss nfet$238
Xpfet$226_0 vdd vdd vosc m1_n8380_274# pfet$226
Xpfet$224_14 vdd m1_n15180_4275# m1_n11782_266# m1_n11916_1270# pfet$224
Xcap_mim$4_0 vss m1_n11296_266# cap_mim$4
Xnfet$238_5 vctrl vss m1_n12754_674# vss nfet$238
Xpfet$226_1 vdd vdd m1_n8380_274# m1_n11916_1270# pfet$226
Xcap_mim$4_1 vss m1_n10810_266# cap_mim$4
Xnfet$238_6 vctrl m1_n16019_266# vss vss nfet$238
Xcap_mim$4_2 vss m1_n10324_266# cap_mim$4
Xnfet$238_7 vctrl vss m1_n15245_186# vss nfet$238
Xpfet$224_0 vdd vdd m1_n12264_2422# m1_n16019_266# pfet$224
Xnfet$238_8 vctrl vss m1_n14765_186# vss nfet$238
Xcap_mim$4_3 vss m1_n11916_1270# cap_mim$4
Xpfet$224_1 vdd vdd m1_n14208_3657# m1_n16019_266# pfet$224
Xnfet$238_9 m1_n10324_266# m1_n13240_368# m1_n9838_266# vss nfet$238
Xcap_mim$4_4 vss m1_n9352_266# cap_mim$4
Xpfet$224_2 vdd vdd m1_n13722_3340# m1_n16019_266# pfet$224
Xcap_mim$4_5 vss m1_n9838_266# cap_mim$4
Xpfet$224_3 vdd m1_n16019_266# vdd m1_n16019_266# pfet$224
Xcap_mim$4_6 vss m1_n11782_266# cap_mim$4
Xpfet$224_4 vdd vdd m1_n13236_3035# m1_n16019_266# pfet$224
Xpfet$224_5 vdd vdd m1_n14693_3963# m1_n16019_266# pfet$224
Xpfet$224_6 vdd vdd m1_n12750_2729# m1_n16019_266# pfet$224
Xpfet$224_7 vdd vdd m1_n15180_4275# m1_n16019_266# pfet$224
Xpfet$224_8 vdd m1_n13236_3035# m1_n9838_266# m1_n10324_266# pfet$224
Xnfet$239_0 vss vss vss vss nfet$239
Xpfet$224_9 vdd m1_n12750_2729# m1_n9352_266# m1_n9838_266# pfet$224
Xnfet$239_1 vss vss vss vss nfet$239
Xnfet$238_10 m1_n9352_266# m1_n12268_985# m1_n11916_1270# vss nfet$238
Xnfet$238_11 m1_n11916_1270# m1_n15245_186# m1_n11782_266# vss nfet$238
Xnfet$238_12 m1_n11782_266# m1_n14765_186# m1_n11296_266# vss nfet$238
Xnfet$238_13 m1_n11296_266# m1_n14283_186# m1_n10810_266# vss nfet$238
Xnfet$238_14 m1_n10810_266# m1_n13794_186# m1_n10324_266# vss nfet$238
Xpfet$225_0 vdd vdd vdd vdd pfet$225
Xnfet$240_0 m1_n8380_274# vss vosc vss nfet$240
Xpfet$225_1 vdd vdd vdd vdd pfet$225
Xnfet$240_1 m1_n11916_1270# vss m1_n8380_274# vss nfet$240
Xnfet$238_0 m1_n9838_266# m1_n12754_674# m1_n9352_266# vss nfet$238
.ends

.subckt top_level_20250912_nosc i_cp_100u div_def div_prc_s8 div_prc_s7 div_prc_s6
+ div_prc_s5 div_prc_s4 div_prc_s3 div_prc_s2 div_prc_s1 div_prc_s0 div_in div_swc_s0
+ div_swc_s1 div_swc_s2 div_swc_s3 div_swc_s4 div_swc_s5 div_swc_s6 div_swc_s7 div_swc_s8
+ lock ref ext_pfd_div ext_pfd_ref ext_pfd_up ext_pfd_down mx_pfd_s1 mx_pfd_s0 down
+ cp_s1 cp_s2 cp_s3 cp_s4 filter_in out filter_out mx_vco_s0 mx_vco_s1 div_rpc_s0
+ div_rsc_s0 div_rsc_s1 div_rpc_s1 div_rsc_s2 div_rpc_s2 div_rsc_s3 div_rsc_s4 div_rsc_s5
+ div_rsc_s6 div_rsc_s7 div_rsc_s8 div_rpc_s3 div_rpc_s4 div_rpc_s5 div_rpc_s6 div_rpc_s7
+ div_rpc_s8 mx_ref_s1 mx_ref_s0 xp_3_1_MUX_1/B_1 up ext_vco_out BIAS_0/200p2 BIAS_0/200p1
+ vdd ext_vco_in BIAS_0/200n div_out vss xp_3_1_MUX_0/B_1
Xasc_drive_buffer_up_0 vss asc_drive_buffer_up_0/out xp_3_1_MUX_2/OUT_1 vdd asc_drive_buffer_up
Xasc_dual_psd_def_20250809_0 vdd vss div_prc_s0 div_prc_s1 div_prc_s2 div_prc_s3 div_prc_s4
+ div_prc_s5 div_prc_s6 div_prc_s7 div_prc_s8 xp_3_1_MUX_4/OUT_1 div_swc_s0 div_swc_s1
+ div_swc_s2 div_swc_s3 div_swc_s4 div_swc_s5 div_swc_s6 div_swc_s7 div_swc_s8 asc_drive_buffer_0/in
+ div_def asc_dual_psd_def_20250809
Xasc_drive_buffer_0 vss asc_drive_buffer_0/in vdd div_in asc_drive_buffer
Xxp_3_1_MUX$1_0 mx_ref_s0 mx_ref_s1 vdd vss xp_3_1_MUX$1_0/OUT_1 xp_3_1_MUX$1_1/C_1
+ xp_3_1_MUX$1_0/B_1 xp_3_1_MUX$1_0/A_1 xp_3_1_MUX$1
Xasc_hysteresis_buffer$2_0 vss ref vdd xp_3_1_MUX$1_0/OUT_1 asc_hysteresis_buffer$2
Xasc_drive_buffer_1 vss xp_3_1_MUX_0/OUT_1 vdd out asc_drive_buffer
Xxp_3_1_MUX$1_1 mx_ref_s0 mx_ref_s1 vdd vss xp_3_1_MUX$1_1/OUT_1 xp_3_1_MUX$1_1/C_1
+ xp_3_1_MUX$1_1/B_1 xp_3_1_MUX$1_1/A_1 xp_3_1_MUX$1
Xasc_drive_buffer_2 vss xp_3_1_MUX_4/OUT_1 vdd div_out asc_drive_buffer
Xasc_drive_buffer_3 vss asc_drive_buffer_3/in vdd lock asc_drive_buffer
Xasc_lock_detector_20250826_0 xp_3_1_MUX_3/OUT_1 vdd xp_3_1_MUX_4/OUT_1 vss asc_drive_buffer_3/in
+ asc_lock_detector_20250826
Xasc_drive_buffer_4 vss xp_3_1_MUX_2/OUT_1 vdd up asc_drive_buffer
Xasc_drive_buffer_5 vss xp_3_1_MUX_5/OUT_1 vdd down asc_drive_buffer
Xasc_drive_buffer_6 vss xp_3_1_MUX_5/OUT_1 vdd asc_drive_buffer_6/out asc_drive_buffer
Xasc_dual_psd_def_20250809$1_0 vdd vss div_rpc_s0 div_rpc_s1 div_rpc_s2 div_rpc_s3
+ div_rpc_s4 div_rpc_s5 div_rpc_s6 div_rpc_s7 div_rpc_s8 xp_3_1_MUX$1_1/B_1 div_rsc_s0
+ div_rsc_s1 div_rsc_s2 div_rsc_s3 div_rsc_s4 div_rsc_s5 div_rsc_s6 div_rsc_s7 div_rsc_s8
+ xp_3_1_MUX$1_0/B_1 vss asc_dual_psd_def_20250809$1
Xasc_drive_buffer$1_0 vss xp_3_1_MUX_0/OUT_1 vdd asc_drive_buffer_0/in asc_drive_buffer$1
Xxp_3_1_MUX_0 mx_vco_s0 mx_vco_s1 vdd vss xp_3_1_MUX_0/OUT_1 xp_3_1_MUX_0/C_1 xp_3_1_MUX_0/B_1
+ ext_vco_out xp_3_1_MUX
Xxp_3_1_MUX_1 mx_vco_s0 mx_vco_s1 vdd vss filter_out xp_3_1_MUX_1/C_1 xp_3_1_MUX_1/B_1
+ ext_vco_in xp_3_1_MUX
Xxp_3_1_MUX_2 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX_2/OUT_1 xp_3_1_MUX_2/C_1 xp_3_1_MUX_2/B_1
+ ext_pfd_up xp_3_1_MUX
Xxp_3_1_MUX_3 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX_3/OUT_1 xp_3_1_MUX_3/C_1 xp_3_1_MUX_3/B_1
+ ext_pfd_ref xp_3_1_MUX
Xxp_3_1_MUX_4 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX_4/OUT_1 xp_3_1_MUX_4/C_1 xp_3_1_MUX_4/B_1
+ ext_pfd_div xp_3_1_MUX
Xxp_programmable_basic_pump_0 asc_drive_buffer_up_0/out vdd cp_s1 cp_s2 cp_s3 cp_s4
+ asc_drive_buffer_6/out filter_in BIAS_0/100n vss xp_programmable_basic_pump
Xxp_3_1_MUX_5 mx_pfd_s0 mx_pfd_s1 vdd vss xp_3_1_MUX_5/OUT_1 xp_3_1_MUX_5/C_1 xp_3_1_MUX_5/B_1
+ ext_pfd_down xp_3_1_MUX
Xasc_hysteresis_buffer$1_0 vss xp_3_1_MUX$1_1/OUT_1 vdd xp_3_1_MUX_3/OUT_1 asc_hysteresis_buffer$1
Xasc_PFD_DFF_20250831_0 vss xp_3_1_MUX_5/C_1 xp_3_1_MUX_2/C_1 vdd xp_3_1_MUX_3/C_1
+ xp_3_1_MUX_4/C_1 asc_PFD_DFF_20250831
XBIAS_0 vdd vss BIAS_0/100n BIAS_0/200n i_cp_100u BIAS_0/200p1 BIAS_0/200p2 BIAS
Xasc_PFD_DFF_20250831_1 vss xp_3_1_MUX_2/B_1 xp_3_1_MUX_5/B_1 vdd xp_3_1_MUX_3/B_1
+ xp_3_1_MUX_4/B_1 asc_PFD_DFF_20250831
XCSRVCO_20250823_0 xp_3_1_MUX_1/C_1 xp_3_1_MUX_0/C_1 vdd vss CSRVCO_20250823
.ends

.subckt pfet$125 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=1.625p ps=6.3u w=2.5u l=0.28u
.ends

.subckt nfet$133 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt pfet$123 a_1054_0# a_734_0# a_254_0# a_894_0# a_348_560# a_828_560# a_988_560#
+ w_n180_n88# a_1214_0# a_414_0# a_n92_0# a_94_0# a_574_0# a_508_560# a_188_560# a_668_560#
+ a_1148_560# a_28_560#
X0 a_1214_0# a_1148_560# a_1054_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_734_0# a_668_560# a_574_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X3 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X4 a_1054_0# a_988_560# a_894_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X5 a_894_0# a_828_560# a_734_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X6 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X7 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt pfet$124 a_254_0# a_348_560# w_n180_n88# a_414_0# a_n92_0# a_94_0# a_574_0#
+ a_508_560# a_188_560# a_28_560#
X0 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$134 a_254_0# a_n84_0# a_94_0# a_190_460# a_30_460# VSUBS
X0 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt nfet$132 a_1054_0# a_734_0# a_510_n132# a_254_0# a_894_0# a_670_n132# a_1214_0#
+ a_830_n132# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132# a_574_0# a_990_n132#
+ a_350_n132# a_1150_n132# VSUBS
X0 a_734_0# a_670_n132# a_574_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X3 a_1054_0# a_990_n132# a_894_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X4 a_894_0# a_830_n132# a_734_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X5 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X6 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X7 a_1214_0# a_1150_n132# a_1054_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt Pcomparator vss vdd out iref inn inp
Xpfet$125_2 vdd vdd vdd vdd pfet$125
Xpfet$125_1 vdd vdd vdd vdd pfet$125
Xnfet$133_1 vss vss vss vss vss vss vss vss vss vss nfet$133
Xnfet$133_0 vss vss vss vss vss vss vss vss vss vss nfet$133
Xpfet$125_3 vdd vdd vdd vdd pfet$125
Xpfet$123_1 out out vdd vdd iref iref iref vdd vdd out vdd out vdd iref iref iref
+ iref iref pfet$123
Xpfet$123_0 out out vdd vdd iref iref iref vdd vdd out vdd out vdd iref iref iref
+ iref iref pfet$123
Xpfet$124_10 vdd iref vdd iref vdd iref vdd iref iref iref pfet$124
Xpfet$124_11 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$124
Xpfet$124_12 m1_2779_n1752# inn vdd m1_3615_n1223# m1_2779_n1752# m1_3615_n1223# m1_2779_n1752#
+ inn inn inn pfet$124
Xpfet$124_13 m1_2779_n1752# inp vdd m1_5539_n2811# m1_2779_n1752# m1_5539_n2811# m1_2779_n1752#
+ inp inp inp pfet$124
Xnfet$134_0 vss vss m1_3615_n1223# m1_3615_n1223# m1_3615_n1223# vss nfet$134
Xnfet$134_1 vss vss m1_5539_n2811# m1_3615_n1223# m1_3615_n1223# vss nfet$134
Xnfet$134_2 vss vss m1_5539_n2811# m1_3615_n1223# m1_3615_n1223# vss nfet$134
Xpfet$124_0 m1_2779_n1752# inp vdd m1_5539_n2811# m1_2779_n1752# m1_5539_n2811# m1_2779_n1752#
+ inp inp inp pfet$124
Xnfet$132_0 out out m1_5539_n2811# vss vss m1_5539_n2811# vss m1_5539_n2811# out m1_5539_n2811#
+ vss out m1_5539_n2811# vss m1_5539_n2811# m1_5539_n2811# m1_5539_n2811# vss nfet$132
Xnfet$134_3 vss vss m1_3615_n1223# m1_3615_n1223# m1_3615_n1223# vss nfet$134
Xpfet$124_1 m1_2779_n1752# m1_2779_n1752# vdd m1_2779_n1752# m1_2779_n1752# m1_2779_n1752#
+ m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# pfet$124
Xpfet$124_2 m1_2779_n1752# inn vdd m1_3615_n1223# m1_2779_n1752# m1_3615_n1223# m1_2779_n1752#
+ inn inn inn pfet$124
Xpfet$124_3 m1_2779_n1752# m1_2779_n1752# vdd m1_2779_n1752# m1_2779_n1752# m1_2779_n1752#
+ m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# m1_2779_n1752# pfet$124
Xpfet$124_4 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$124
Xpfet$124_6 vdd iref vdd iref vdd iref vdd iref iref iref pfet$124
Xpfet$124_5 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$124
Xpfet$124_7 vdd iref vdd iref vdd iref vdd iref iref iref pfet$124
Xpfet$124_8 vdd iref vdd iref vdd iref vdd iref iref iref pfet$124
Xpfet$124_9 vdd iref vdd m1_2779_n1752# vdd m1_2779_n1752# vdd iref iref iref pfet$124
Xpfet$125_0 vdd vdd vdd vdd pfet$125
.ends

.subckt nfet$128 a_254_0# a_n84_0# a_94_0# a_190_460# a_30_460# VSUBS
X0 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt nfet$131 a_n84_0# a_94_0# a_30_460# VSUBS
X0 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$121 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
.ends

.subckt nfet$129 a_1054_0# a_734_0# a_254_0# a_350_460# a_830_460# a_894_0# a_990_460#
+ a_1214_0# a_414_0# a_n84_0# a_94_0# a_510_460# a_190_460# a_574_0# a_670_460# a_1150_460#
+ a_30_460# VSUBS
X0 a_734_0# a_670_460# a_574_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_574_0# a_510_460# a_414_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X3 a_1054_0# a_990_460# a_894_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X4 a_894_0# a_830_460# a_734_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X5 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X6 a_414_0# a_350_460# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X7 a_1214_0# a_1150_460# a_1054_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt pfet$122 a_254_0# a_348_560# w_n180_n88# a_414_0# a_n92_0# a_94_0# a_574_0#
+ a_508_560# a_188_560# a_28_560#
X0 a_254_0# a_188_560# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_560# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_560# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_560# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$130 a_254_0# a_350_460# a_414_0# a_n84_0# a_94_0# a_510_460# a_190_460#
+ a_574_0# a_30_460# VSUBS
X0 a_254_0# a_190_460# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_460# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_460# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt pfet$120 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_348_n136# a_414_0#
+ a_n92_0# a_94_0# a_574_0# a_508_n136#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_n136# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_n136# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt Ncomparator vss vdd out inn inp iref
Xnfet$128_3 m1_506_n191# m1_506_n191# m1_1242_549# inn inn vss nfet$128
Xnfet$131_0 vss vss vss vss nfet$131
Xnfet$131_1 vss vss vss vss nfet$131
Xpfet$121_0 vdd vdd vdd vdd vdd vdd pfet$121
Xpfet$121_1 vdd vdd vdd vdd vdd vdd pfet$121
Xpfet$121_2 vdd vdd vdd vdd vdd vdd pfet$121
Xpfet$121_3 vdd vdd vdd vdd vdd vdd pfet$121
Xnfet$129_0 out out vss iref iref vss iref vss out vss out iref iref vss iref iref
+ iref vss nfet$129
Xpfet$122_0 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$122
Xpfet$122_1 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$122
Xnfet$130_0 vss iref m1_506_n191# vss m1_506_n191# iref iref vss iref vss nfet$130
Xpfet$122_2 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$122
Xnfet$130_1 vss iref iref vss iref iref iref vss iref vss nfet$130
Xpfet$120_0 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_570_1653# vdd m1_570_1653#
+ vdd m1_1242_549# pfet$120
Xpfet$122_3 vdd m1_570_1653# vdd out vdd out vdd m1_570_1653# m1_570_1653# m1_570_1653#
+ pfet$122
Xnfet$130_3 m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191#
+ m1_506_n191# m1_506_n191# m1_506_n191# vss nfet$130
Xnfet$130_2 m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191# m1_506_n191#
+ m1_506_n191# m1_506_n191# m1_506_n191# vss nfet$130
Xpfet$120_1 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_1242_549# vdd m1_1242_549#
+ vdd m1_1242_549# pfet$120
Xnfet$130_4 vss iref iref vss iref iref iref vss iref vss nfet$130
Xpfet$120_3 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_1242_549# vdd m1_1242_549#
+ vdd m1_1242_549# pfet$120
Xpfet$120_2 m1_1242_549# vdd m1_1242_549# vdd m1_1242_549# m1_570_1653# vdd m1_570_1653#
+ vdd m1_1242_549# pfet$120
Xnfet$130_5 vss iref m1_506_n191# vss m1_506_n191# iref iref vss iref vss nfet$130
Xnfet$128_1 m1_506_n191# m1_506_n191# m1_1242_549# inn inn vss nfet$128
Xnfet$128_0 m1_506_n191# m1_506_n191# m1_570_1653# inp inp vss nfet$128
Xnfet$128_2 m1_506_n191# m1_506_n191# m1_570_1653# inp inp vss nfet$128
.ends

.subckt nfet$13 a_n84_0# a_94_0# a_30_160# VSUBS
X0 a_94_0# a_30_160# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=0.28u
.ends

.subckt pfet$12 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt SRLATCH vdd vss q qb s r
Xnfet$13_0 vss qb r vss nfet$13
Xnfet$13_1 vss qb q vss nfet$13
Xpfet$12_0 r vdd m1_818_875# qb pfet$12
Xnfet$13_2 q vss s vss nfet$13
Xpfet$12_1 q vdd vdd m1_818_875# pfet$12
Xnfet$13_3 q vss qb vss nfet$13
Xpfet$12_2 s vdd m1_50_875# vdd pfet$12
Xpfet$12_3 qb vdd q m1_50_875# pfet$12
.ends

.subckt ppolyf_u_resistor$2 a_n376_0# a_4200_0# a_n132_0#
X0 a_n132_0# a_4200_0# a_n376_0# ppolyf_u r_width=1u r_length=21u
.ends

.subckt pfet$128 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt nfet$136 a_30_n132# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$126 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=2.6p pd=9.3u as=2.6p ps=9.3u w=4u l=0.28u
.ends

.subckt pfet$127 a_28_460# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_460# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt nfet$135 a_n84_0# a_94_0# a_30_460# VSUBS
X0 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt SCHMITT VDD VSS IN OUT
Xnfet$136_0 OUT m1_592_402# VDD VSS nfet$136
Xpfet$126_0 IN VDD m1_596_1544# OUT pfet$126
Xpfet$126_1 IN VDD VDD m1_596_1544# pfet$126
Xpfet$127_0 OUT VDD m1_596_1544# VSS pfet$127
Xnfet$135_0 m1_592_402# OUT IN VSS nfet$135
Xnfet$135_1 VSS m1_592_402# IN VSS nfet$135
.ends

.subckt cap_mim$3 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=60u c_length=100u
.ends

.subckt nfet$137 a_30_260# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_260# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.28u
.ends

.subckt pfet$118 a_750_0# a_546_0# a_446_n60# a_242_n60# w_n180_n88# a_38_n60# a_n92_0#
+ a_342_0# a_138_0# a_650_n60#
X0 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X2 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.5u
.ends

.subckt nfet$126 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.5u
.ends

.subckt nfet$122 a_750_0# a_546_0# a_446_n132# a_n84_0# a_650_n132# a_38_n132# a_342_0#
+ a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.5u
X1 a_546_0# a_446_n132# a_342_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.5u
X2 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.5u
X3 a_750_0# a_650_n132# a_546_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.5u
.ends

.subckt pfet$116 a_28_460# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_460# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt nfet$124 a_750_0# a_546_0# a_446_n132# a_n84_0# a_650_n132# a_38_n132# a_342_0#
+ a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_546_0# a_446_n132# a_342_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.26p ps=1.52u w=1u l=0.5u
X2 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
X3 a_750_0# a_650_n132# a_546_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt pfet$114 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# w_n180_n88# a_1262_n60# a_38_n60# a_n92_0# a_1058_n60# a_854_n60# a_342_0#
+ a_138_0# a_650_n60# a_1362_0#
X0 a_1362_0# a_1262_n60# a_1158_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X1 a_954_0# a_854_n60# a_750_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X2 a_1566_0# a_1466_n60# a_1362_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.5u
X3 a_342_0# a_242_n60# a_138_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X4 a_546_0# a_446_n60# a_342_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X5 a_1158_0# a_1058_n60# a_954_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
X6 a_138_0# a_38_n60# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.5u
X7 a_750_0# a_650_n60# a_546_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.5u
.ends

.subckt cap_mim$2 m4_n120_n120# m4_0_0#
X0 m4_0_0# m4_n120_n120# cap_mim_2f0_m4m5_noshield c_width=50u c_length=100u
.ends

.subckt nfet$119 a_254_0# a_30_n132# a_n84_0# a_94_0# a_190_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$112 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_348_n136# a_414_0#
+ a_n92_0# a_94_0# a_574_0# a_508_n136#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_574_0# a_508_n136# a_414_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X3 a_414_0# a_348_n136# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$120 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt pfet$113 a_28_n136# a_254_0# a_188_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
.ends

.subckt OTAforChargePump$1 vdd vss out iref inn inp
Xnfet$119_0 vss m1_116_n1334# vss out m1_116_n1334# vss nfet$119
Xnfet$119_1 vss m1_116_n1334# vss m1_116_n1334# m1_116_n1334# vss nfet$119
Xnfet$119_2 vss m1_116_n1334# vss m1_116_n1334# m1_116_n1334# vss nfet$119
Xnfet$119_3 vss m1_116_n1334# vss out m1_116_n1334# vss nfet$119
Xpfet$112_0 inn m1_n400_n914# inn vdd inn out m1_n400_n914# out m1_n400_n914# inn
+ pfet$112
Xpfet$112_1 inp m1_n400_n914# inp vdd inp m1_116_n1334# m1_n400_n914# m1_116_n1334#
+ m1_n400_n914# inp pfet$112
Xnfet$120_0 vss vss vss vss vss vss vss vss vss vss nfet$120
Xpfet$112_2 iref vdd iref vdd iref iref vdd iref vdd iref pfet$112
Xnfet$120_1 vss vss vss vss vss vss vss vss vss vss nfet$120
Xpfet$112_3 iref vdd iref vdd iref m1_n400_n914# vdd m1_n400_n914# vdd iref pfet$112
Xpfet$112_4 iref vdd iref vdd iref m1_n400_n914# vdd m1_n400_n914# vdd iref pfet$112
Xpfet$112_6 iref vdd iref vdd iref iref vdd iref vdd iref pfet$112
Xpfet$112_5 iref vdd iref vdd iref iref vdd iref vdd iref pfet$112
Xpfet$112_7 iref vdd iref vdd iref m1_n400_n914# vdd m1_n400_n914# vdd iref pfet$112
Xpfet$112_8 inp m1_n400_n914# inp vdd inp m1_116_n1334# m1_n400_n914# m1_116_n1334#
+ m1_n400_n914# inp pfet$112
Xpfet$112_9 inn m1_n400_n914# inn vdd inn out m1_n400_n914# out m1_n400_n914# inn
+ pfet$112
Xpfet$113_0 m1_n400_n914# m1_n400_n914# m1_n400_n914# vdd m1_n400_n914# m1_n400_n914#
+ pfet$113
Xpfet$113_2 vdd vdd vdd vdd vdd vdd pfet$113
Xpfet$113_1 m1_n400_n914# m1_n400_n914# m1_n400_n914# vdd m1_n400_n914# m1_n400_n914#
+ pfet$113
Xpfet$113_3 vdd vdd vdd vdd vdd vdd pfet$113
Xpfet$113_4 vdd vdd vdd vdd vdd vdd pfet$113
Xpfet$113_5 vdd vdd vdd vdd vdd vdd pfet$113
Xpfet$112_10 iref vdd iref vdd iref iref vdd iref vdd iref pfet$112
Xpfet$112_11 iref vdd iref vdd iref m1_n400_n914# vdd m1_n400_n914# vdd iref pfet$112
.ends

.subckt pfet$119 a_1054_0# a_734_0# a_828_n136# a_28_n136# a_254_0# a_894_0# a_188_n136#
+ a_988_n136# w_n180_n88# a_348_n136# a_1214_0# a_1148_n136# a_414_0# a_n92_0# a_94_0#
+ a_574_0# a_508_n136# a_668_n136#
X0 a_1214_0# a_1148_n136# a_1054_0# w_n180_n88# pfet_03v3 ad=1.625p pd=6.3u as=0.65p ps=3.02u w=2.5u l=0.28u
X1 a_734_0# a_668_n136# a_574_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X2 a_254_0# a_188_n136# a_94_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X3 a_574_0# a_508_n136# a_414_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X4 a_1054_0# a_988_n136# a_894_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X5 a_894_0# a_828_n136# a_734_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
X6 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=1.625p ps=6.3u w=2.5u l=0.28u
X7 a_414_0# a_348_n136# a_254_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.02u as=0.65p ps=3.02u w=2.5u l=0.28u
.ends

.subckt nfet$127 a_510_n132# a_254_0# a_414_0# a_30_n132# a_n84_0# a_94_0# a_190_n132#
+ a_574_0# a_350_n132# VSUBS
X0 a_254_0# a_190_n132# a_94_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
X1 a_574_0# a_510_n132# a_414_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=0.52p ps=2.52u w=2u l=0.28u
X2 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=1.22p ps=5.22u w=2u l=0.28u
X3 a_414_0# a_350_n132# a_254_0# VSUBS nfet_03v3 ad=0.52p pd=2.52u as=0.52p ps=2.52u w=2u l=0.28u
.ends

.subckt pfet$117 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$125 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$115 w_n180_n88# a_n92_0# a_342_0# a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=0.8125p pd=3.8u as=0.325p ps=1.77u w=1.25u l=0.5u
X1 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.325p pd=1.77u as=0.8125p ps=3.8u w=1.25u l=0.5u
.ends

.subckt nfet$123 a_n84_0# a_38_n132# a_342_0# a_138_0# a_242_n132# VSUBS
X0 a_342_0# a_242_n132# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n132# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt nfet$121 a_30_n132# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt ppolyf_u_resistor$1 a_4000_0# a_n376_0# a_n132_0#
X0 a_n132_0# a_4000_0# a_n376_0# ppolyf_u r_width=1u r_length=20u
.ends

.subckt PCP1248X vdd vss s3 s2 s1 s0 vin iref200u out up down
Xpfet$118_11 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$118
Xpfet$118_0 m1_n47_11059# m1_n47_11059# m1_n47_11059# m1_n47_11059# vdd m1_n47_11059#
+ m1_n47_11059# m1_n47_11059# m1_n47_11059# m1_n47_11059# pfet$118
Xpfet$118_1 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$118
Xnfet$126_0 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$126
Xpfet$118_2 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$118
Xnfet$122_30 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$122
Xnfet$126_1 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$126
Xpfet$118_3 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$118
Xnfet$126_2 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$126
Xnfet$122_20 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$122
Xpfet$116_0 s0 vdd m1_1641_5849# vdd pfet$116
Xnfet$122_31 m1_n47_11059# m1_14015_1164# m1_9963_14448# m1_n47_11059# m1_9963_14448#
+ m1_9963_14448# m1_n47_11059# m1_14015_1164# m1_9963_14448# vss nfet$122
Xpfet$118_4 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$118
Xnfet$122_21 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$122
Xnfet$126_3 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$126
Xnfet$122_32 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$122
Xnfet$122_10 m1_13543_n1758# m1_15911_n1318# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15911_n1318# m1_9963_14448# vss nfet$122
Xnfet$124_0 vss m1_9475_12045# OTAforChargePump$1_0/out vss OTAforChargePump$1_0/out
+ OTAforChargePump$1_0/out vss m1_9475_12045# OTAforChargePump$1_0/out vss nfet$124
Xpfet$116_1 s3 vdd m1_n1771_4009# vdd pfet$116
Xnfet$126_4 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ vss nfet$126
Xnfet$124_1 vss m1_n1751_n2187# OTAforChargePump$1_0/out vss OTAforChargePump$1_0/out
+ OTAforChargePump$1_0/out vss m1_n1751_n2187# OTAforChargePump$1_0/out vss nfet$124
Xnfet$122_22 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$122
Xnfet$122_33 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$122
Xpfet$116_2 m1_n1311_12403# vdd m1_n47_11059# m1_n91_6229# pfet$116
Xnfet$122_11 m1_13543_n1758# m1_15039_784# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15039_784# m1_9963_14448# vss nfet$122
Xpfet$118_5 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$118
Xnfet$122_34 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$122
Xnfet$122_23 vss m1_15039_784# m1_15009_5932# vss m1_15009_5932# m1_15009_5932# vss
+ m1_15039_784# m1_15009_5932# vss nfet$122
Xpfet$118_6 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$118
Xnfet$126_5 m1_n47_11059# m1_n47_11059# m1_n47_11059# m1_n47_11059# m1_n47_11059#
+ vss nfet$126
Xnfet$122_12 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$122
Xnfet$124_2 vss m1_9475_12045# OTAforChargePump$1_0/out vss OTAforChargePump$1_0/out
+ OTAforChargePump$1_0/out vss m1_9475_12045# OTAforChargePump$1_0/out vss nfet$124
Xpfet$116_3 m1_n2083_12403# vdd m1_n47_11059# m1_1137_12199# pfet$116
Xpfet$114_0 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$114
Xnfet$126_6 vss vss vss vss vss vss nfet$126
Xnfet$124_3 vss m1_n1751_n2187# OTAforChargePump$1_0/out vss OTAforChargePump$1_0/out
+ OTAforChargePump$1_0/out vss m1_n1751_n2187# OTAforChargePump$1_0/out vss nfet$124
Xnfet$122_24 vss vss vss vss vss vss vss vss vss vss nfet$122
Xnfet$122_35 vss m1_14015_1164# OTAforChargePump$1_0/out vss OTAforChargePump$1_0/out
+ OTAforChargePump$1_0/out vss m1_14015_1164# OTAforChargePump$1_0/out vss nfet$122
Xpfet$118_7 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$118
Xpfet$116_4 m1_n2855_12403# vdd m1_n47_11059# m1_n1771_4009# pfet$116
Xnfet$122_13 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$122
Xcap_mim$2_0 m1_n1751_n2187# vdd cap_mim$2
Xpfet$114_1 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$114
Xnfet$122_0 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$122
Xnfet$126_7 vss vss vss vss vss vss nfet$126
Xpfet$118_8 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# pfet$118
Xcap_mim$2_1 vss m1_9963_14448# cap_mim$2
Xnfet$122_36 OTAforChargePump$1_0/inp m1_9475_12045# m1_9963_14448# OTAforChargePump$1_0/inp
+ m1_9963_14448# m1_9963_14448# OTAforChargePump$1_0/inp m1_9475_12045# m1_9963_14448#
+ vss nfet$122
Xnfet$122_25 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$122
Xpfet$116_5 s1 vdd m1_n91_6229# vdd pfet$116
Xnfet$122_1 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$122
Xnfet$122_14 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$122
Xpfet$114_2 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$114
Xnfet$126_8 vss vss vss vss vss vss nfet$126
Xnfet$122_26 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$122
Xnfet$122_15 vss vss vss vss vss vss vss vss vss vss nfet$122
Xpfet$118_9 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$118
Xpfet$116_6 s2 vdd m1_1137_12199# vdd pfet$116
Xcap_mim$2_2 vss OTAforChargePump$1_0/out cap_mim$2
Xnfet$122_2 m1_13543_n1758# m1_14167_n938# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_14167_n938# m1_9963_14448# vss nfet$122
Xpfet$114_3 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$114
Xnfet$126_9 vss vss vss vss vss vss nfet$126
Xnfet$122_27 vss m1_15911_n1318# m1_15881_3450# vss m1_15881_3450# m1_15881_3450#
+ vss m1_15911_n1318# m1_15881_3450# vss nfet$122
Xnfet$122_16 vss m1_16783_404# m1_16753_5552# vss m1_16753_5552# m1_16753_5552# vss
+ m1_16783_404# m1_16753_5552# vss nfet$122
Xpfet$116_7 m1_n539_12403# vdd m1_n47_11059# m1_1641_5849# pfet$116
Xnfet$122_3 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# vss nfet$122
Xpfet$116_10 m1_n2083_12403# vdd OTAforChargePump$1_0/out m1_15881_3450# pfet$116
Xpfet$114_4 m1_n2925_n36# m1_n2925_n36# m1_n25_493# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n25_493# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36#
+ m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n25_493# m1_n1751_n2187# m1_n25_493#
+ pfet$114
Xnfet$122_28 vss m1_15911_n1318# m1_15881_3450# vss m1_15881_3450# m1_15881_3450#
+ vss m1_15911_n1318# m1_15881_3450# vss nfet$122
Xnfet$122_17 vss m1_15039_784# m1_15009_5932# vss m1_15009_5932# m1_15009_5932# vss
+ m1_15039_784# m1_15009_5932# vss nfet$122
Xpfet$116_8 m1_n539_12403# vdd OTAforChargePump$1_0/out m1_16753_5552# pfet$116
Xpfet$114_5 m1_n47_11059# m1_n47_11059# m1_6759_7857# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n47_11059# m1_6759_7857# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n47_11059# m1_n1751_n2187# m1_n1751_n2187# m1_n47_11059# m1_6759_7857# m1_n1751_n2187#
+ m1_6759_7857# pfet$114
Xnfet$122_4 m1_13543_n1758# m1_15039_784# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15039_784# m1_9963_14448# vss nfet$122
Xpfet$116_11 m1_n2855_12403# vdd OTAforChargePump$1_0/out m1_14137_3830# pfet$116
Xpfet$116_9 m1_n1311_12403# vdd OTAforChargePump$1_0/out m1_15009_5932# pfet$116
Xnfet$122_29 vss m1_14167_n938# m1_14137_3830# vss m1_14137_3830# m1_14137_3830# vss
+ m1_14167_n938# m1_14137_3830# vss nfet$122
Xnfet$122_18 vss m1_15911_n1318# m1_15881_3450# vss m1_15881_3450# m1_15881_3450#
+ vss m1_15911_n1318# m1_15881_3450# vss nfet$122
Xpfet$114_6 vdd vdd m1_6759_7857# m1_n47_11059# m1_n47_11059# vdd m1_6759_7857# m1_n47_11059#
+ vdd m1_n47_11059# m1_n47_11059# vdd m1_n47_11059# m1_n47_11059# vdd m1_6759_7857#
+ m1_n47_11059# m1_6759_7857# pfet$114
XOTAforChargePump$1_0 vdd vss OTAforChargePump$1_0/out iref200u vin OTAforChargePump$1_0/inp
+ OTAforChargePump$1
Xnfet$122_5 m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758#
+ m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# m1_13543_n1758# vss nfet$122
Xnfet$122_19 vss m1_15911_n1318# m1_15881_3450# vss m1_15881_3450# m1_15881_3450#
+ vss m1_15911_n1318# m1_15881_3450# vss nfet$122
Xpfet$114_7 vdd vdd m1_n25_493# m1_n91_6229# m1_n91_6229# vdd m1_n25_493# m1_n91_6229#
+ vdd m1_n91_6229# m1_n91_6229# vdd m1_n91_6229# m1_n91_6229# vdd m1_n25_493# m1_n91_6229#
+ m1_n25_493# pfet$114
Xnfet$122_6 m1_13543_n1758# m1_16783_404# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_16783_404# m1_9963_14448# vss nfet$122
Xnfet$122_7 m1_13543_n1758# m1_15911_n1318# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15911_n1318# m1_9963_14448# vss nfet$122
Xpfet$114_8 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$114
Xnfet$122_8 m1_13543_n1758# m1_15911_n1318# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15911_n1318# m1_9963_14448# vss nfet$122
Xpfet$114_9 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$114
Xpfet$119_0 m1_n2925_n36# m1_n2925_n36# up up out out up up vdd up out up m1_n2925_n36#
+ out m1_n2925_n36# out up up pfet$119
Xnfet$122_9 m1_13543_n1758# m1_15911_n1318# m1_9963_14448# m1_13543_n1758# m1_9963_14448#
+ m1_9963_14448# m1_13543_n1758# m1_15911_n1318# m1_9963_14448# vss nfet$122
Xnfet$126_10 vss vss vss vss vss vss nfet$126
Xnfet$127_0 down out m1_13543_n1758# down out m1_13543_n1758# down out down vss nfet$127
Xnfet$126_11 vss vss vss vss vss vss nfet$126
Xpfet$117_0 vdd vdd m1_n2855_12403# s3 pfet$117
Xpfet$114_30 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ pfet$114
Xpfet$117_1 vdd vdd m1_n2083_12403# s2 pfet$117
Xnfet$125_0 s3 vss m1_n2855_12403# vss nfet$125
Xpfet$114_31 m1_n2925_n36# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187#
+ m1_1671_n1319# pfet$114
Xpfet$114_20 m1_n2925_n36# m1_n2925_n36# m1_1671_873# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_873# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36#
+ m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_873# m1_n1751_n2187# m1_1671_873#
+ pfet$114
Xnfet$125_1 s2 vss m1_n2083_12403# vss nfet$125
Xpfet$117_2 vdd vdd m1_n539_12403# s0 pfet$117
Xpfet$114_10 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$114
Xpfet$114_32 m1_n2925_n36# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187#
+ m1_1671_n1319# pfet$114
Xpfet$114_21 vdd vdd m1_1671_873# m1_1641_5849# m1_1641_5849# vdd m1_1671_873# m1_1641_5849#
+ vdd m1_1641_5849# m1_1641_5849# vdd m1_1641_5849# m1_1641_5849# vdd m1_1671_873#
+ m1_1641_5849# m1_1671_873# pfet$114
Xpfet$117_3 vdd vdd m1_n1311_12403# s1 pfet$117
Xnfet$125_2 s1 vss m1_n1311_12403# vss nfet$125
Xpfet$115_0 vdd vdd vdd vdd vdd vdd pfet$115
Xpfet$114_11 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$114
Xpfet$114_22 vdd vdd m1_1671_n1319# m1_1137_12199# m1_1137_12199# vdd m1_1671_n1319#
+ m1_1137_12199# vdd m1_1137_12199# m1_1137_12199# vdd m1_1137_12199# m1_1137_12199#
+ vdd m1_1671_n1319# m1_1137_12199# m1_1671_n1319# pfet$114
Xpfet$114_33 vdd vdd m1_1671_n1319# m1_1137_12199# m1_1137_12199# vdd m1_1671_n1319#
+ m1_1137_12199# vdd m1_1137_12199# m1_1137_12199# vdd m1_1137_12199# m1_1137_12199#
+ vdd m1_1671_n1319# m1_1137_12199# m1_1671_n1319# pfet$114
Xnfet$125_3 s0 vss m1_n539_12403# vss nfet$125
Xpfet$115_1 vdd vdd vdd m1_n1751_n2187# m1_n1751_n2187# m1_n1751_n2187# pfet$115
Xnfet$123_0 vss vss vss vss vss vss nfet$123
Xpfet$114_12 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$114
Xpfet$114_23 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$114
Xpfet$114_34 vdd vdd m1_1671_n1319# m1_1137_12199# m1_1137_12199# vdd m1_1671_n1319#
+ m1_1137_12199# vdd m1_1137_12199# m1_1137_12199# vdd m1_1137_12199# m1_1137_12199#
+ vdd m1_1671_n1319# m1_1137_12199# m1_1671_n1319# pfet$114
Xnfet$123_1 vss vss vss vss vss vss nfet$123
Xpfet$115_2 vdd vdd vdd m1_9963_14448# m1_n1751_n2187# m1_n1751_n2187# pfet$115
Xpfet$114_13 m1_n2925_n36# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187#
+ m1_1671_n1319# pfet$114
Xpfet$114_24 vdd vdd m1_n25_493# m1_n91_6229# m1_n91_6229# vdd m1_n25_493# m1_n91_6229#
+ vdd m1_n91_6229# m1_n91_6229# vdd m1_n91_6229# m1_n91_6229# vdd m1_n25_493# m1_n91_6229#
+ m1_n25_493# pfet$114
Xpfet$114_35 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ pfet$114
Xpfet$115_3 vdd vdd vdd m1_n1751_n2187# m1_n1751_n2187# m1_n1751_n2187# pfet$115
Xnfet$123_2 vss m1_9963_14448# vss m1_9963_14448# m1_9963_14448# vss nfet$123
Xpfet$114_14 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$114
Xpfet$114_25 vdd vdd m1_1671_n1319# m1_1137_12199# m1_1137_12199# vdd m1_1671_n1319#
+ m1_1137_12199# vdd m1_1137_12199# m1_1137_12199# vdd m1_1137_12199# m1_1137_12199#
+ vdd m1_1671_n1319# m1_1137_12199# m1_1671_n1319# pfet$114
Xpfet$115_4 vdd vdd vdd m1_9963_14448# m1_n1751_n2187# m1_n1751_n2187# pfet$115
Xnfet$121_0 s0 m1_n47_11059# m1_1641_5849# vss nfet$121
Xpfet$114_15 m1_n2925_n36# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_1671_n1319# m1_n1751_n2187#
+ m1_1671_n1319# pfet$114
Xpfet$114_26 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$114
Xnfet$121_10 m1_n2855_12403# m1_14137_3830# vss vss nfet$121
Xpfet$115_5 vdd vdd vdd vdd vdd vdd pfet$115
Xnfet$121_1 s1 m1_n47_11059# m1_n91_6229# vss nfet$121
Xpfet$114_16 m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# vdd m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36# m1_n2925_n36#
+ pfet$114
Xpfet$114_27 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$114
Xnfet$121_11 s3 OTAforChargePump$1_0/out m1_14137_3830# vss nfet$121
Xpfet$114_17 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$114
Xpfet$114_28 vdd vdd m1_n1721_n939# m1_n1771_4009# m1_n1771_4009# vdd m1_n1721_n939#
+ m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009# vdd m1_n1771_4009# m1_n1771_4009#
+ vdd m1_n1721_n939# m1_n1771_4009# m1_n1721_n939# pfet$114
Xnfet$121_2 s3 m1_n47_11059# m1_n1771_4009# vss nfet$121
Xppolyf_u_resistor$1_0 m1_3630_13790# vss m1_n502_13390# ppolyf_u_resistor$1
Xnfet$121_3 s2 m1_n47_11059# m1_1137_12199# vss nfet$121
Xpfet$114_18 m1_n2925_n36# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n1721_n939# m1_n1751_n2187#
+ m1_n1721_n939# pfet$114
Xpfet$114_29 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd
+ pfet$114
Xppolyf_u_resistor$1_1 OTAforChargePump$1_0/inp vss m1_n502_13390# ppolyf_u_resistor$1
Xnfet$121_4 m1_n539_12403# m1_16753_5552# vss vss nfet$121
Xpfet$114_19 m1_n2925_n36# m1_n2925_n36# m1_n25_493# m1_n1751_n2187# m1_n1751_n2187#
+ m1_n2925_n36# m1_n25_493# m1_n1751_n2187# vdd m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36#
+ m1_n1751_n2187# m1_n1751_n2187# m1_n2925_n36# m1_n25_493# m1_n1751_n2187# m1_n25_493#
+ pfet$114
Xppolyf_u_resistor$1_2 m1_3630_14590# vss m1_n502_14190# ppolyf_u_resistor$1
Xnfet$121_5 s0 OTAforChargePump$1_0/out m1_16753_5552# vss nfet$121
Xppolyf_u_resistor$1_3 m1_3630_13790# vss m1_n502_14190# ppolyf_u_resistor$1
Xnfet$121_6 m1_n1311_12403# m1_15009_5932# vss vss nfet$121
Xppolyf_u_resistor$1_4 m1_3630_14590# vss m1_n502_14990# ppolyf_u_resistor$1
Xnfet$121_7 s1 OTAforChargePump$1_0/out m1_15009_5932# vss nfet$121
Xppolyf_u_resistor$1_5 vdd vss m1_n502_14990# ppolyf_u_resistor$1
Xnfet$121_8 m1_n2083_12403# m1_15881_3450# vss vss nfet$121
Xpfet$118_10 vdd vdd vdd vdd vdd vdd vdd vdd vdd vdd pfet$118
Xnfet$121_9 s2 OTAforChargePump$1_0/out m1_15881_3450# vss nfet$121
.ends

.subckt VCOfinal vdd s3 iref200 fout foutb irefn irefp s1 s2 a_11641_n18839# s0 vin
+ vss
XPcomparator_0 vss vdd SRLATCH_0/r irefp PCP1248X_0/out Pcomparator_0/inp Pcomparator
XNcomparator_0 vss vdd SRLATCH_0/s Ncomparator_0/inn PCP1248X_0/out irefn Ncomparator
XSRLATCH_0 vdd vss SRLATCH_0/q SRLATCH_0/qb SRLATCH_0/s SRLATCH_0/r SRLATCH
Xppolyf_u_resistor$2_0 vss vss Pcomparator_0/inp ppolyf_u_resistor$2
Xppolyf_u_resistor$2_1 vss m1_13996_n13334# Ncomparator_0/inn ppolyf_u_resistor$2
Xpfet$128_0 SRLATCH_0/q vdd vdd PCP1248X_0/up pfet$128
Xppolyf_u_resistor$2_2 vss m1_13996_n13334# Pcomparator_0/inp ppolyf_u_resistor$2
Xpfet$128_1 SCHMITT_0/OUT vdd vdd foutb pfet$128
Xppolyf_u_resistor$2_3 vss vdd Ncomparator_0/inn ppolyf_u_resistor$2
Xpfet$128_2 SCHMITT_1/OUT vdd vdd fout pfet$128
XSCHMITT_0 vdd vss SRLATCH_0/qb SCHMITT_0/OUT SCHMITT
XSCHMITT_1 vdd vss SRLATCH_0/q SCHMITT_1/OUT SCHMITT
Xcap_mim$3_0 vss PCP1248X_0/out cap_mim$3
Xnfet$137_0 SRLATCH_0/q vss PCP1248X_0/up vss nfet$137
Xnfet$137_1 SCHMITT_0/OUT vss foutb vss nfet$137
XPCP1248X_0 vdd vss s3 s2 s1 s0 vin iref200 PCP1248X_0/out PCP1248X_0/up SRLATCH_0/qb
+ PCP1248X
Xnfet$137_2 SCHMITT_1/OUT vss fout vss nfet$137
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__and2_1$2 A1 A2 VDD VSS Z VNW VPW
X0 VDD A2 a_36_201# VNW pfet_05v0 ad=0.5054p pd=2.57u as=0.2132p ps=1.34u w=0.82u l=0.5u
X1 a_244_201# A1 a_36_201# VPW nfet_05v0 ad=0.1056p pd=0.98u as=0.2904p ps=2.2u w=0.66u l=0.6u
X2 Z a_36_201# VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.3894p ps=2.06u w=1.32u l=0.6u
X3 Z a_36_201# VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.5054p ps=2.57u w=1.83u l=0.5u
X4 VSS A2 a_244_201# VPW nfet_05v0 ad=0.3894p pd=2.06u as=0.1056p ps=0.98u w=0.66u l=0.6u
X5 a_36_201# A1 VDD VNW pfet_05v0 ad=0.2132p pd=1.34u as=0.3608p ps=2.52u w=0.82u l=0.5u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__or2_1$2 A1 A2 VDD VSS Z VNW VPW
X0 a_255_756# A1 a_67_756# VNW pfet_05v0 ad=0.2379p pd=1.435u as=0.4026p ps=2.71u w=0.915u l=0.5u
X1 VSS A2 a_67_756# VPW nfet_05v0 ad=0.3828p pd=2.08u as=0.1716p ps=1.18u w=0.66u l=0.6u
X2 VDD A2 a_255_756# VNW pfet_05v0 ad=0.57645p pd=2.69u as=0.2379p ps=1.435u w=0.915u l=0.5u
X3 Z a_67_756# VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.3828p ps=2.08u w=1.32u l=0.6u
X4 Z a_67_756# VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.57645p ps=2.69u w=1.83u l=0.5u
X5 a_67_756# A1 VSS VPW nfet_05v0 ad=0.1716p pd=1.18u as=0.2904p ps=2.2u w=0.66u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__inv_1$2 I VDD VSS ZN VNW VPW
X0 ZN I VDD VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X1 ZN I VSS VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
.ends

.subckt gf180mcu_fd_sc_mcu9t5v0__latq_1$3 D E Q VDD VSS VNW VPW
X0 VSS a_1020_652# Q VPW nfet_05v0 ad=0.5808p pd=3.52u as=0.5808p ps=3.52u w=1.32u l=0.6u
X1 a_504_110# a_36_92# VDD VNW pfet_05v0 ad=0.44p pd=2.88u as=0.476p ps=2.18u w=1u l=0.5u
X2 VDD a_1020_652# Q VNW pfet_05v0 ad=0.8052p pd=4.54u as=0.8052p ps=4.54u w=1.83u l=0.5u
X3 a_1264_107# a_36_92# a_1020_652# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.182p ps=1.22u w=0.7u l=0.6u
X4 VSS E a_36_92# VPW nfet_05v0 ad=0.263p pd=1.49u as=0.3476p ps=2.46u w=0.79u l=0.6u
X5 VSS a_1364_532# a_1264_107# VPW nfet_05v0 ad=0.2054p pd=1.31u as=0.263p ps=1.49u w=0.79u l=0.6u
X6 VDD E a_36_92# VNW pfet_05v0 ad=0.476p pd=2.18u as=0.6072p ps=3.64u w=1.38u l=0.5u
X7 VDD a_1364_532# a_1224_652# VNW pfet_05v0 ad=0.3588p pd=1.9u as=0.426p ps=2.08u w=1.38u l=0.5u
X8 a_872_652# D VDD VNW pfet_05v0 ad=0.12p pd=1.24u as=0.44p ps=2.88u w=1u l=0.5u
X9 a_1364_532# a_1020_652# VDD VNW pfet_05v0 ad=0.6072p pd=3.64u as=0.3588p ps=1.9u w=1.38u l=0.5u
X10 a_1020_652# a_504_110# a_872_107# VPW nfet_05v0 ad=0.182p pd=1.22u as=83.99999f ps=0.94u w=0.7u l=0.6u
X11 a_872_107# D VSS VPW nfet_05v0 ad=83.99999f pd=0.94u as=0.308p ps=2.28u w=0.7u l=0.6u
X12 a_1020_652# a_36_92# a_872_652# VNW pfet_05v0 ad=0.26p pd=1.52u as=0.12p ps=1.24u w=1u l=0.5u
X13 a_504_110# a_36_92# VSS VPW nfet_05v0 ad=0.308p pd=2.28u as=0.263p ps=1.49u w=0.7u l=0.6u
X14 a_1364_532# a_1020_652# VSS VPW nfet_05v0 ad=0.3476p pd=2.46u as=0.2054p ps=1.31u w=0.79u l=0.6u
X15 a_1224_652# a_504_110# a_1020_652# VNW pfet_05v0 ad=0.426p pd=2.08u as=0.26p ps=1.52u w=1u l=0.5u
.ends

.subckt DFF_2phase_1$2 VDDd PHI_1 D Q PHI_2 VSSd
Xgf180mcu_fd_sc_mcu9t5v0__latq_1$3_0 gf180mcu_fd_sc_mcu9t5v0__latq_1$3_1/Q PHI_2 Q
+ VDDd VSSd VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1$3
Xgf180mcu_fd_sc_mcu9t5v0__latq_1$3_1 D PHI_1 gf180mcu_fd_sc_mcu9t5v0__latq_1$3_1/Q
+ VDDd VSSd VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__latq_1$3
.ends

.subckt Register_unitcell$1 out d q en default phi1 phi2 VSSd VDDd
Xgf180mcu_fd_sc_mcu9t5v0__and2_1$2_0 gf180mcu_fd_sc_mcu9t5v0__inv_1$2_0/ZN default
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1$2_0/A1 VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1$2
Xgf180mcu_fd_sc_mcu9t5v0__and2_1$2_1 q en VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1$2_0/A2
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__and2_1$2
Xgf180mcu_fd_sc_mcu9t5v0__or2_1$2_0 gf180mcu_fd_sc_mcu9t5v0__or2_1$2_0/A1 gf180mcu_fd_sc_mcu9t5v0__or2_1$2_0/A2
+ VDDd VSSd out VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__or2_1$2
Xgf180mcu_fd_sc_mcu9t5v0__inv_1$2_0 en VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1$2_0/ZN
+ VDDd VSSd gf180mcu_fd_sc_mcu9t5v0__inv_1$2
XDFF_2phase_1$2_0 VDDd phi1 d q phi2 VSSd DFF_2phase_1$2
.ends

.subckt SRegister_10 out[1] out[2] out[3] out[8] d default10 default9 default8 default7
+ default6 default5 default4 default3 default2 default1 out[9] out[6] out[4] out[10]
+ out[7] phi2 out[5] en phi1 q VSSd VDDd
XRegister_unitcell$1_0 out[2] Register_unitcell$1_6/q Register_unitcell$1_7/d en default2
+ phi1 phi2 VSSd VDDd Register_unitcell$1
XRegister_unitcell$1_1 out[6] Register_unitcell$1_9/q Register_unitcell$1_2/d en default6
+ phi1 phi2 VSSd VDDd Register_unitcell$1
XRegister_unitcell$1_2 out[7] Register_unitcell$1_2/d Register_unitcell$1_3/d en default7
+ phi1 phi2 VSSd VDDd Register_unitcell$1
XRegister_unitcell$1_3 out[8] Register_unitcell$1_3/d Register_unitcell$1_4/d en default8
+ phi1 phi2 VSSd VDDd Register_unitcell$1
XRegister_unitcell$1_4 out[9] Register_unitcell$1_4/d Register_unitcell$1_5/d en default9
+ phi1 phi2 VSSd VDDd Register_unitcell$1
XRegister_unitcell$1_5 out[10] Register_unitcell$1_5/d q en default10 phi1 phi2 VSSd
+ VDDd Register_unitcell$1
XRegister_unitcell$1_7 out[3] Register_unitcell$1_7/d Register_unitcell$1_8/d en default3
+ phi1 phi2 VSSd VDDd Register_unitcell$1
XRegister_unitcell$1_6 out[1] d Register_unitcell$1_6/q en default1 phi1 phi2 VSSd
+ VDDd Register_unitcell$1
XRegister_unitcell$1_8 out[4] Register_unitcell$1_8/d Register_unitcell$1_9/d en default4
+ phi1 phi2 VSSd VDDd Register_unitcell$1
XRegister_unitcell$1_9 out[5] Register_unitcell$1_9/d Register_unitcell$1_9/q en default5
+ phi1 phi2 VSSd VDDd Register_unitcell$1
.ends

.subckt pfet$139 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$147 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$137 a_838_0# w_n180_n88# a_n92_0# a_38_n136#
X0 a_838_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=4u
.ends

.subckt nfet$145 a_38_n60# a_n84_0# a_438_0# VSUBS
X0 a_438_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=2u
.ends

.subckt nfet$148 a_242_n60# a_38_n60# a_n84_0# a_342_0# a_138_0# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.26p ps=1.52u w=1u l=0.5u
X1 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.26p pd=1.52u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$138 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$146 a_838_0# a_38_n60# a_n84_0# VSUBS
X0 a_838_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.305p pd=2.22u as=0.305p ps=2.22u w=0.5u l=4u
.ends

.subckt pfet$136 w_n180_n88# a_n92_0# a_438_0# a_38_n136#
X0 a_438_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=0.65p pd=3.3u as=0.65p ps=3.3u w=1u l=2u
.ends

.subckt qw_NOLclk VDDd VSSd PHI_1 PHI_2 CLK
Xpfet$139_0 VDDd m1_11601_71# VDDd m1_11379_n171# pfet$139
Xnfet$147_0 m1_11601_71# VSSd PHI_1 VSSd nfet$147
Xpfet$139_1 VDDd VDDd m1_11601_71# m1_12351_431# pfet$139
Xpfet$139_2 VDDd m1_11601_2380# VDDd m1_11161_409# pfet$139
Xnfet$147_1 m1_11161_409# VSSd m1_11379_n171# VSSd nfet$147
Xpfet$139_3 VDDd VDDd m1_11601_2380# m1_12351_2064# pfet$139
Xnfet$147_2 m1_11601_2380# VSSd PHI_2 VSSd nfet$147
Xnfet$147_3 CLK VSSd m1_11161_409# VSSd nfet$147
Xpfet$137_0 m1_12351_2064# VDDd VDDd m1_15103_233# pfet$137
Xpfet$137_2 m1_12351_431# VDDd VDDd m1_15103_1818# pfet$137
Xnfet$145_1 PHI_2 VSSd m1_13930_1818# VSSd nfet$145
Xnfet$145_0 PHI_1 VSSd m1_13930_233# VSSd nfet$145
Xpfet$137_1 m1_15103_233# VDDd VDDd m1_13930_233# pfet$137
Xpfet$137_3 m1_15103_1818# VDDd VDDd m1_13930_1818# pfet$137
Xnfet$148_0 m1_12351_431# m1_12351_431# m1_11601_71# m1_11601_71# m1_11837_749# VSSd
+ nfet$148
Xnfet$148_1 m1_11379_n171# m1_11379_n171# VSSd VSSd m1_11837_749# VSSd nfet$148
Xnfet$148_2 m1_12351_2064# m1_12351_2064# m1_11601_2380# m1_11601_2380# m1_11837_1708#
+ VSSd nfet$148
Xpfet$138_0 VDDd VDDd PHI_1 m1_11601_71# pfet$138
Xnfet$148_3 m1_11161_409# m1_11161_409# VSSd VSSd m1_11837_1708# VSSd nfet$148
Xnfet$146_0 m1_12351_2064# m1_15103_233# VSSd VSSd nfet$146
Xpfet$138_1 VDDd VDDd m1_11379_n171# m1_11161_409# pfet$138
Xpfet$138_2 VDDd VDDd PHI_2 m1_11601_2380# pfet$138
Xnfet$146_1 m1_15103_233# m1_13930_233# VSSd VSSd nfet$146
Xpfet$138_3 VDDd VDDd m1_11161_409# CLK pfet$138
Xnfet$146_2 m1_12351_431# m1_15103_1818# VSSd VSSd nfet$146
Xpfet$136_0 VDDd VDDd m1_13930_233# PHI_1 pfet$136
Xpfet$136_1 VDDd VDDd m1_13930_1818# PHI_2 pfet$136
Xnfet$146_3 m1_15103_1818# m1_13930_1818# VSSd VSSd nfet$146
.ends

.subckt pfet$135 a_28_460# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_460# a_n92_0# w_n180_n88# pfet_03v3 ad=1.3p pd=5.3u as=1.3p ps=5.3u w=2u l=0.28u
.ends

.subckt nfet$143 a_n84_0# a_94_0# a_30_460# VSUBS
X0 a_94_0# a_30_460# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt nfet$144 a_30_n132# a_n84_0# a_94_0# VSUBS
X0 a_94_0# a_30_n132# a_n84_0# VSUBS nfet_03v3 ad=1.22p pd=5.22u as=1.22p ps=5.22u w=2u l=0.28u
.ends

.subckt pfet$134 a_28_n136# w_n180_n88# a_n92_0# a_94_0#
X0 a_94_0# a_28_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=2.6p pd=9.3u as=2.6p ps=9.3u w=4u l=0.28u
.ends

.subckt SCHMITT$1 VDD VSS IN OUT
Xpfet$135_0 OUT VDD m1_596_1544# VSS pfet$135
Xnfet$143_0 m1_592_402# OUT IN VSS nfet$143
Xnfet$143_1 VSS m1_592_402# IN VSS nfet$143
Xnfet$144_0 OUT m1_592_402# VDD VSS nfet$144
Xpfet$134_0 IN VDD m1_596_1544# OUT pfet$134
Xpfet$134_1 IN VDD VDD m1_596_1544# pfet$134
.ends

.subckt pfet$130 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$138 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$133 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$141 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$131 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$139 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$129 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$142 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$132 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$140 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_hysteresis_buffer vss in vdd out
Xpfet$130_0 vdd vdd m1_884_42# m1_348_648# pfet$130
Xnfet$138_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$138
Xpfet$133_0 vdd vdd m1_884_42# m1_1156_42# pfet$133
Xnfet$141_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$141
Xpfet$131_0 vdd vdd m1_348_648# in pfet$131
Xnfet$139_0 m1_348_648# vss m1_884_42# vss nfet$139
Xpfet$129_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd
+ m1_884_42# m1_884_42# pfet$129
Xnfet$142_0 m1_1156_42# vss m1_884_42# vss nfet$142
Xpfet$132_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$132
Xnfet$140_0 in vss m1_348_648# vss nfet$140
.ends

.subckt scan_chain VDDd ENd DATAd CLKd out[1] out[2] out[3] out[4] out[5] out[6] out[7]
+ out[8] out[9] out[10] out[20] out[19] out[18] out[17] out[16] out[15] out[14] out[13]
+ out[12] out[11] out[21] out[22] out[23] out[24] out[25] out[26] out[27] out[28]
+ out[29] out[30] out[40] out[39] out[38] out[37] out[36] out[35] out[34] out[33]
+ out[32] out[31] out[41] out[42] out[43] out[44] out[45] out[46] out[47] out[48]
+ out[49] out[50] VSSd
XSRegister_10_1 out[11] out[12] out[13] out[18] SRegister_10_4/q VSSd VSSd VSSd VSSd
+ VSSd VSSd VSSd VSSd VSSd VSSd out[19] out[16] out[14] out[20] out[17] qw_NOLclk_0/PHI_2
+ out[15] SRegister_10_4/en qw_NOLclk_0/PHI_1 SRegister_10_3/d VSSd VDDd SRegister_10
XSRegister_10_2 out[41] out[42] out[43] out[48] SRegister_10_2/d VSSd VSSd VSSd VSSd
+ VDDd VSSd VSSd VDDd VDDd VSSd out[49] out[46] out[44] out[50] out[47] qw_NOLclk_0/PHI_2
+ out[45] SRegister_10_4/en qw_NOLclk_0/PHI_1 SRegister_10_2/q VSSd VDDd SRegister_10
Xqw_NOLclk_0 VDDd VSSd qw_NOLclk_0/PHI_1 qw_NOLclk_0/PHI_2 qw_NOLclk_0/CLK qw_NOLclk
XSRegister_10_3 out[21] out[22] out[23] out[28] SRegister_10_3/d VSSd VSSd VSSd VSSd
+ VSSd VSSd VSSd VSSd VSSd VSSd out[29] out[26] out[24] out[30] out[27] qw_NOLclk_0/PHI_2
+ out[25] SRegister_10_4/en qw_NOLclk_0/PHI_1 SRegister_10_3/q VSSd VDDd SRegister_10
XSCHMITT$1_0 VDDd VSSd SCHMITT$1_0/IN qw_NOLclk_0/CLK SCHMITT$1
XSRegister_10_4 out[1] out[2] out[3] out[8] SRegister_10_4/d VSSd VSSd VSSd VSSd VDDd
+ VSSd VSSd VSSd VSSd VSSd out[9] out[6] out[4] out[10] out[7] qw_NOLclk_0/PHI_2 out[5]
+ SRegister_10_4/en qw_NOLclk_0/PHI_1 SRegister_10_4/q VSSd VDDd SRegister_10
Xasc_hysteresis_buffer_0 VSSd CLKd VDDd SCHMITT$1_0/IN asc_hysteresis_buffer
Xasc_hysteresis_buffer_1 VSSd ENd VDDd SRegister_10_4/en asc_hysteresis_buffer
Xasc_hysteresis_buffer_2 VSSd DATAd VDDd SRegister_10_4/d asc_hysteresis_buffer
XSRegister_10_0 out[31] out[32] out[33] out[38] SRegister_10_3/q VSSd VSSd VDDd VSSd
+ VSSd VDDd VDDd VSSd VSSd VSSd out[39] out[36] out[34] out[40] out[37] qw_NOLclk_0/PHI_2
+ out[35] SRegister_10_4/en qw_NOLclk_0/PHI_1 SRegister_10_2/d VSSd VDDd SRegister_10
.ends

.subckt nfet$29 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt pfet$28 a_1158_0# a_750_0# a_1058_n136# a_546_0# a_1262_n136# a_1566_0# a_954_0#
+ w_n180_n88# a_854_n136# a_n92_0# a_446_n136# a_650_n136# a_342_0# a_1466_n136# a_138_0#
+ a_38_n136# a_1362_0# a_242_n136#
X0 a_1362_0# a_1262_n136# a_1158_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_954_0# a_854_n136# a_750_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_1566_0# a_1466_n136# a_1362_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
X3 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X4 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X5 a_1158_0# a_1058_n136# a_954_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X6 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X7 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$27 a_750_0# a_546_0# a_446_n60# a_242_n60# a_38_n60# a_n84_0# a_342_0#
+ a_138_0# a_650_n60# VSUBS
X0 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X3 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$26 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=7.8p ps=25.3u w=12u l=0.5u
.ends

.subckt nfet$30 a_1158_0# a_750_0# a_546_0# a_446_n60# a_242_n60# a_1566_0# a_954_0#
+ a_1466_n60# a_1262_n60# a_38_n60# a_n84_0# a_1058_n60# a_854_n60# a_342_0# a_138_0#
+ a_650_n60# a_1362_0# VSUBS
X0 a_954_0# a_854_n60# a_750_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X1 a_1566_0# a_1466_n60# a_1362_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=1.04p ps=4.52u w=4u l=0.5u
X2 a_342_0# a_242_n60# a_138_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X3 a_546_0# a_446_n60# a_342_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X4 a_1158_0# a_1058_n60# a_954_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X5 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=2.44p ps=9.22u w=4u l=0.5u
X6 a_750_0# a_650_n60# a_546_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
X7 a_1362_0# a_1262_n60# a_1158_0# VSUBS nfet_03v3 ad=1.04p pd=4.52u as=1.04p ps=4.52u w=4u l=0.5u
.ends

.subckt pfet$29 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt nfet$28 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=2.44p pd=9.22u as=2.44p ps=9.22u w=4u l=0.5u
.ends

.subckt pfet$27 w_n180_n88# a_n92_0# a_138_0# a_38_n136#
X0 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=1.95p pd=7.3u as=1.95p ps=7.3u w=3u l=0.5u
.ends

.subckt pfet$25 a_750_0# a_546_0# w_n180_n88# a_n92_0# a_446_n136# a_650_n136# a_342_0#
+ a_138_0# a_38_n136# a_242_n136#
X0 a_342_0# a_242_n136# a_138_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X1 a_546_0# a_446_n136# a_342_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=3.12p ps=12.52u w=12u l=0.5u
X2 a_138_0# a_38_n136# a_n92_0# w_n180_n88# pfet_03v3 ad=3.12p pd=12.52u as=7.8p ps=25.3u w=12u l=0.5u
X3 a_750_0# a_650_n136# a_546_0# w_n180_n88# pfet_03v3 ad=7.8p pd=25.3u as=3.12p ps=12.52u w=12u l=0.5u
.ends

.subckt nfet$31 a_38_n60# a_n84_0# a_138_0# VSUBS
X0 a_138_0# a_38_n60# a_n84_0# VSUBS nfet_03v3 ad=0.61p pd=3.22u as=0.61p ps=3.22u w=1u l=0.5u
.ends

.subckt asc_hysteresis_buffer$3 vss vdd out in
Xnfet$29_0 in vss m1_348_648# vss nfet$29
Xpfet$28_0 out out m1_1156_42# vdd m1_1156_42# out vdd vdd m1_1156_42# out m1_1156_42#
+ m1_1156_42# out m1_1156_42# vdd m1_1156_42# vdd m1_1156_42# pfet$28
Xnfet$27_0 m1_1156_42# vss m1_884_42# m1_884_42# m1_884_42# m1_1156_42# m1_1156_42#
+ vss m1_884_42# vss nfet$27
Xpfet$26_0 vdd vdd m1_884_42# m1_348_648# pfet$26
Xnfet$30_0 out out vss m1_1156_42# m1_1156_42# out vss m1_1156_42# m1_1156_42# m1_1156_42#
+ out m1_1156_42# m1_1156_42# out vss m1_1156_42# vss vss nfet$30
Xpfet$29_0 vdd vdd m1_884_42# m1_1156_42# pfet$29
Xnfet$28_0 m1_348_648# vss m1_884_42# vss nfet$28
Xpfet$27_0 vdd vdd m1_348_648# in pfet$27
Xpfet$25_0 m1_1156_42# vdd vdd m1_1156_42# m1_884_42# m1_884_42# m1_1156_42# vdd m1_884_42#
+ m1_884_42# pfet$25
Xnfet$31_0 m1_1156_42# vss m1_884_42# vss nfet$31
.ends

.subckt top_level_20250919_sc VDDd VSSd en clk data div_def ref ext_pfd_div ext_pfd_ref
+ ext_pfd_down ext_pfd_up i_cp_100u up down lock filter_in filter_out ext_vco_in ext_vco_out
+ out div_in div_out
Xtop_level_20250912_nosc_0 i_cp_100u asc_hysteresis_buffer$3_0/out scan_chain_0/out[42]
+ scan_chain_0/out[43] scan_chain_0/out[44] scan_chain_0/out[45] scan_chain_0/out[46]
+ scan_chain_0/out[47] scan_chain_0/out[48] scan_chain_0/out[49] scan_chain_0/out[50]
+ div_in scan_chain_0/out[41] scan_chain_0/out[40] scan_chain_0/out[39] scan_chain_0/out[38]
+ scan_chain_0/out[37] scan_chain_0/out[36] scan_chain_0/out[35] scan_chain_0/out[34]
+ scan_chain_0/out[33] lock ref ext_pfd_div ext_pfd_ref ext_pfd_up ext_pfd_down scan_chain_0/out[1]
+ scan_chain_0/out[2] down scan_chain_0/out[6] scan_chain_0/out[5] scan_chain_0/out[4]
+ scan_chain_0/out[3] filter_in out filter_out scan_chain_0/out[32] scan_chain_0/out[31]
+ scan_chain_0/out[26] scan_chain_0/out[17] scan_chain_0/out[16] scan_chain_0/out[25]
+ scan_chain_0/out[15] scan_chain_0/out[24] scan_chain_0/out[14] scan_chain_0/out[13]
+ scan_chain_0/out[12] scan_chain_0/out[11] scan_chain_0/out[10] scan_chain_0/out[9]
+ scan_chain_0/out[23] scan_chain_0/out[22] scan_chain_0/out[21] scan_chain_0/out[20]
+ scan_chain_0/out[19] scan_chain_0/out[18] scan_chain_0/out[7] scan_chain_0/out[8]
+ VCOfinal_0/vin up ext_vco_out VCOfinal_0/irefp VCOfinal_0/iref200 VDDd ext_vco_in
+ VCOfinal_0/irefn div_out VSSd VCOfinal_0/fout top_level_20250912_nosc
XVCOfinal_0 VDDd VCOfinal_0/s3 VCOfinal_0/iref200 VCOfinal_0/fout VCOfinal_0/foutb
+ VCOfinal_0/irefn VCOfinal_0/irefp VCOfinal_0/s1 VCOfinal_0/s2 VSSd VCOfinal_0/s0
+ VCOfinal_0/vin VSSd VCOfinal
Xscan_chain_0 VDDd en data clk scan_chain_0/out[1] scan_chain_0/out[2] scan_chain_0/out[3]
+ scan_chain_0/out[4] scan_chain_0/out[5] scan_chain_0/out[6] scan_chain_0/out[7]
+ scan_chain_0/out[8] scan_chain_0/out[9] scan_chain_0/out[10] scan_chain_0/out[20]
+ scan_chain_0/out[19] scan_chain_0/out[18] scan_chain_0/out[17] scan_chain_0/out[16]
+ scan_chain_0/out[15] scan_chain_0/out[14] scan_chain_0/out[13] scan_chain_0/out[12]
+ scan_chain_0/out[11] scan_chain_0/out[21] scan_chain_0/out[22] scan_chain_0/out[23]
+ scan_chain_0/out[24] scan_chain_0/out[25] scan_chain_0/out[26] VCOfinal_0/s0 VCOfinal_0/s1
+ VCOfinal_0/s2 VCOfinal_0/s3 scan_chain_0/out[40] scan_chain_0/out[39] scan_chain_0/out[38]
+ scan_chain_0/out[37] scan_chain_0/out[36] scan_chain_0/out[35] scan_chain_0/out[34]
+ scan_chain_0/out[33] scan_chain_0/out[32] scan_chain_0/out[31] scan_chain_0/out[41]
+ scan_chain_0/out[42] scan_chain_0/out[43] scan_chain_0/out[44] scan_chain_0/out[45]
+ scan_chain_0/out[46] scan_chain_0/out[47] scan_chain_0/out[48] scan_chain_0/out[49]
+ scan_chain_0/out[50] VSSd scan_chain
Xasc_hysteresis_buffer$3_0 VSSd VDDd asc_hysteresis_buffer$3_0/out div_def asc_hysteresis_buffer$3
.ends

