** sch_path: /foss/designs/libs/core_analog/asc_drive_buffer/asc_drive_buffer.sch
.subckt asc_drive_buffer in vss out vdd
*.PININFO in:B out:B vss:B vdd:B
XM1 net1 in vdd vdd pfet_03v3 L=0.5u W=3.0u nf=1 m=1
XM2 net1 in vss vss nfet_03v3 L=0.5u W=1.0u nf=1 m=1
XM3 net2 net1 vdd vdd pfet_03v3 L=0.5u W=12.0u nf=1 m=1
XM4 net2 net1 vss vss nfet_03v3 L=0.5u W=4.0u nf=1 m=1
XM5 net3 net2 vdd vdd pfet_03v3 L=0.5u W=48.0u nf=4 m=1
XM6 net3 net2 vss vss nfet_03v3 L=0.5u W=16.0u nf=4 m=1
XM7 out net3 vdd vdd pfet_03v3 L=0.5u W=96.0u nf=8 m=1
XM8 out net3 vss vss nfet_03v3 L=0.5u W=32.0u nf=8 m=1
.ends
