** sch_path: /foss/designs/libs/core_analog/asc_XNOR/asc_XNOR.sch
.subckt asc_XNOR VDD VSS OUT A B
*.PININFO VDD:B VSS:B B:B A:B OUT:B
M1 OUT A net1 VSS nfet_03v3 L=0.5u W=2u nf=2 m=1
M2 OUT B net3 VDD pfet_03v3 L=0.5u W=6u nf=2 m=1
M3 net1 Bb VSS VSS nfet_03v3 L=0.5u W=2u nf=2 m=1
M4 net3 A VDD VDD pfet_03v3 L=0.5u W=6u nf=2 m=1
M5 OUT Ab net2 VSS nfet_03v3 L=0.5u W=2u nf=2 m=1
M6 OUT Bb net4 VDD pfet_03v3 L=0.5u W=6u nf=2 m=1
M7 net2 B VSS VSS nfet_03v3 L=0.5u W=2u nf=2 m=1
M8 net4 Ab VDD VDD pfet_03v3 L=0.5u W=6u nf=2 m=1
x1 A VDD Ab VSS inv1u05u
x2 B VDD Bb VSS inv1u05u
.ends

* expanding   symbol:  libs/core_analog/inv1u05u/inv1u05u.sym # of pins=4
** sym_path: /foss/designs/libs/core_analog/inv1u05u/inv1u05u.sym
** sch_path: /foss/designs/libs/core_analog/inv1u05u/inv1u05u.sch
.subckt inv1u05u in vdd out vss
*.PININFO in:B out:B vss:B vdd:B
M1 out in vdd vdd pfet_03v3 L=0.5u W=3.0u nf=1 m=1
M2 out in vss vss nfet_03v3 L=0.5u W=1.0u nf=1 m=1
.ends

